

`timescale 1 ns / 1 ps
module kernel0_kernel0 (
  input s_axi_control_AWVALID,
  output s_axi_control_AWREADY,
  input [6-1:0] s_axi_control_AWADDR,
  input s_axi_control_WVALID,
  output s_axi_control_WREADY,
  input [32-1:0] s_axi_control_WDATA,
  input [32/8-1:0] s_axi_control_WSTRB,
  input s_axi_control_ARVALID,
  output s_axi_control_ARREADY,
  input [6-1:0] s_axi_control_ARADDR,
  output s_axi_control_RVALID,
  input s_axi_control_RREADY,
  output [32-1:0] s_axi_control_RDATA,
  output [1:0] s_axi_control_RRESP,
  output s_axi_control_BVALID,
  input s_axi_control_BREADY,
  output [1:0] s_axi_control_BRESP,
  input ap_clk,
  input ap_rst_n,
  output interrupt,
  output m_axi_gmem_cin_AWVALID,
  input m_axi_gmem_cin_AWREADY,
  output [64-1:0] m_axi_gmem_cin_AWADDR,
  output [1-1:0] m_axi_gmem_cin_AWID,
  output [7:0] m_axi_gmem_cin_AWLEN,
  output [2:0] m_axi_gmem_cin_AWSIZE,
  output [1:0] m_axi_gmem_cin_AWBURST,
  output [1:0] m_axi_gmem_cin_AWLOCK,
  output [3:0] m_axi_gmem_cin_AWCACHE,
  output [2:0] m_axi_gmem_cin_AWPROT,
  output [3:0] m_axi_gmem_cin_AWQOS,
  output [3:0] m_axi_gmem_cin_AWREGION,
  output [1-1:0] m_axi_gmem_cin_AWUSER,
  output m_axi_gmem_cin_WVALID,
  input m_axi_gmem_cin_WREADY,
  output [512-1:0] m_axi_gmem_cin_WDATA,
  output [512/8-1:0] m_axi_gmem_cin_WSTRB,
  output m_axi_gmem_cin_WLAST,
  output [1-1:0] m_axi_gmem_cin_WID,
  output [1-1:0] m_axi_gmem_cin_WUSER,
  output m_axi_gmem_cin_ARVALID,
  input m_axi_gmem_cin_ARREADY,
  output [64-1:0] m_axi_gmem_cin_ARADDR,
  output [1-1:0] m_axi_gmem_cin_ARID,
  output [7:0] m_axi_gmem_cin_ARLEN,
  output [2:0] m_axi_gmem_cin_ARSIZE,
  output [1:0] m_axi_gmem_cin_ARBURST,
  output [1:0] m_axi_gmem_cin_ARLOCK,
  output [3:0] m_axi_gmem_cin_ARCACHE,
  output [2:0] m_axi_gmem_cin_ARPROT,
  output [3:0] m_axi_gmem_cin_ARQOS,
  output [3:0] m_axi_gmem_cin_ARREGION,
  output [1-1:0] m_axi_gmem_cin_ARUSER,
  input m_axi_gmem_cin_RVALID,
  output m_axi_gmem_cin_RREADY,
  input [512-1:0] m_axi_gmem_cin_RDATA,
  input m_axi_gmem_cin_RLAST,
  input [1-1:0] m_axi_gmem_cin_RID,
  input [1-1:0] m_axi_gmem_cin_RUSER,
  input [1:0] m_axi_gmem_cin_RRESP,
  input m_axi_gmem_cin_BVALID,
  output m_axi_gmem_cin_BREADY,
  input [1:0] m_axi_gmem_cin_BRESP,
  input [1-1:0] m_axi_gmem_cin_BID,
  input [1-1:0] m_axi_gmem_cin_BUSER,
  output m_axi_gmem_cout_AWVALID,
  input m_axi_gmem_cout_AWREADY,
  output [64-1:0] m_axi_gmem_cout_AWADDR,
  output [1-1:0] m_axi_gmem_cout_AWID,
  output [7:0] m_axi_gmem_cout_AWLEN,
  output [2:0] m_axi_gmem_cout_AWSIZE,
  output [1:0] m_axi_gmem_cout_AWBURST,
  output [1:0] m_axi_gmem_cout_AWLOCK,
  output [3:0] m_axi_gmem_cout_AWCACHE,
  output [2:0] m_axi_gmem_cout_AWPROT,
  output [3:0] m_axi_gmem_cout_AWQOS,
  output [3:0] m_axi_gmem_cout_AWREGION,
  output [1-1:0] m_axi_gmem_cout_AWUSER,
  output m_axi_gmem_cout_WVALID,
  input m_axi_gmem_cout_WREADY,
  output [512-1:0] m_axi_gmem_cout_WDATA,
  output [512/8-1:0] m_axi_gmem_cout_WSTRB,
  output m_axi_gmem_cout_WLAST,
  output [1-1:0] m_axi_gmem_cout_WID,
  output [1-1:0] m_axi_gmem_cout_WUSER,
  output m_axi_gmem_cout_ARVALID,
  input m_axi_gmem_cout_ARREADY,
  output [64-1:0] m_axi_gmem_cout_ARADDR,
  output [1-1:0] m_axi_gmem_cout_ARID,
  output [7:0] m_axi_gmem_cout_ARLEN,
  output [2:0] m_axi_gmem_cout_ARSIZE,
  output [1:0] m_axi_gmem_cout_ARBURST,
  output [1:0] m_axi_gmem_cout_ARLOCK,
  output [3:0] m_axi_gmem_cout_ARCACHE,
  output [2:0] m_axi_gmem_cout_ARPROT,
  output [3:0] m_axi_gmem_cout_ARQOS,
  output [3:0] m_axi_gmem_cout_ARREGION,
  output [1-1:0] m_axi_gmem_cout_ARUSER,
  input m_axi_gmem_cout_RVALID,
  output m_axi_gmem_cout_RREADY,
  input [512-1:0] m_axi_gmem_cout_RDATA,
  input m_axi_gmem_cout_RLAST,
  input [1-1:0] m_axi_gmem_cout_RID,
  input [1-1:0] m_axi_gmem_cout_RUSER,
  input [1:0] m_axi_gmem_cout_RRESP,
  input m_axi_gmem_cout_BVALID,
  output m_axi_gmem_cout_BREADY,
  input [1:0] m_axi_gmem_cout_BRESP,
  input [1-1:0] m_axi_gmem_cout_BID,
  input [1-1:0] m_axi_gmem_cout_BUSER,
  output m_axi_gmem_w_AWVALID,
  input m_axi_gmem_w_AWREADY,
  output [64-1:0] m_axi_gmem_w_AWADDR,
  output [1-1:0] m_axi_gmem_w_AWID,
  output [7:0] m_axi_gmem_w_AWLEN,
  output [2:0] m_axi_gmem_w_AWSIZE,
  output [1:0] m_axi_gmem_w_AWBURST,
  output [1:0] m_axi_gmem_w_AWLOCK,
  output [3:0] m_axi_gmem_w_AWCACHE,
  output [2:0] m_axi_gmem_w_AWPROT,
  output [3:0] m_axi_gmem_w_AWQOS,
  output [3:0] m_axi_gmem_w_AWREGION,
  output [1-1:0] m_axi_gmem_w_AWUSER,
  output m_axi_gmem_w_WVALID,
  input m_axi_gmem_w_WREADY,
  output [512-1:0] m_axi_gmem_w_WDATA,
  output [512/8-1:0] m_axi_gmem_w_WSTRB,
  output m_axi_gmem_w_WLAST,
  output [1-1:0] m_axi_gmem_w_WID,
  output [1-1:0] m_axi_gmem_w_WUSER,
  output m_axi_gmem_w_ARVALID,
  input m_axi_gmem_w_ARREADY,
  output [64-1:0] m_axi_gmem_w_ARADDR,
  output [1-1:0] m_axi_gmem_w_ARID,
  output [7:0] m_axi_gmem_w_ARLEN,
  output [2:0] m_axi_gmem_w_ARSIZE,
  output [1:0] m_axi_gmem_w_ARBURST,
  output [1:0] m_axi_gmem_w_ARLOCK,
  output [3:0] m_axi_gmem_w_ARCACHE,
  output [2:0] m_axi_gmem_w_ARPROT,
  output [3:0] m_axi_gmem_w_ARQOS,
  output [3:0] m_axi_gmem_w_ARREGION,
  output [1-1:0] m_axi_gmem_w_ARUSER,
  input m_axi_gmem_w_RVALID,
  output m_axi_gmem_w_RREADY,
  input [512-1:0] m_axi_gmem_w_RDATA,
  input m_axi_gmem_w_RLAST,
  input [1-1:0] m_axi_gmem_w_RID,
  input [1-1:0] m_axi_gmem_w_RUSER,
  input [1:0] m_axi_gmem_w_RRESP,
  input m_axi_gmem_w_BVALID,
  output m_axi_gmem_w_BREADY,
  input [1:0] m_axi_gmem_w_BRESP,
  input [1-1:0] m_axi_gmem_w_BID,
  input [1-1:0] m_axi_gmem_w_BUSER
);

  parameter C_S_AXI_CONTROL_DATA_WIDTH = 32;
  parameter C_S_AXI_CONTROL_ADDR_WIDTH = 6;
  parameter C_S_AXI_DATA_WIDTH = 32;
  parameter C_S_AXI_ADDR_WIDTH = 32;
  parameter C_M_AXI_GMEM_CIN_ID_WIDTH = 1;
  parameter C_M_AXI_GMEM_CIN_ADDR_WIDTH = 64;
  parameter C_M_AXI_GMEM_CIN_DATA_WIDTH = 512;
  parameter C_M_AXI_GMEM_CIN_AWUSER_WIDTH = 1;
  parameter C_M_AXI_GMEM_CIN_ARUSER_WIDTH = 1;
  parameter C_M_AXI_GMEM_CIN_WUSER_WIDTH = 1;
  parameter C_M_AXI_GMEM_CIN_RUSER_WIDTH = 1;
  parameter C_M_AXI_GMEM_CIN_BUSER_WIDTH = 1;
  parameter C_M_AXI_GMEM_CIN_USER_VALUE = 0;
  parameter C_M_AXI_GMEM_CIN_PROT_VALUE = 0;
  parameter C_M_AXI_GMEM_CIN_CACHE_VALUE = 3;
  parameter C_M_AXI_ID_WIDTH = 1;
  parameter C_M_AXI_ADDR_WIDTH = 64;
  parameter C_M_AXI_DATA_WIDTH = 32;
  parameter C_M_AXI_AWUSER_WIDTH = 1;
  parameter C_M_AXI_ARUSER_WIDTH = 1;
  parameter C_M_AXI_WUSER_WIDTH = 1;
  parameter C_M_AXI_RUSER_WIDTH = 1;
  parameter C_M_AXI_BUSER_WIDTH = 1;
  parameter C_M_AXI_GMEM_COUT_ID_WIDTH = 1;
  parameter C_M_AXI_GMEM_COUT_ADDR_WIDTH = 64;
  parameter C_M_AXI_GMEM_COUT_DATA_WIDTH = 512;
  parameter C_M_AXI_GMEM_COUT_AWUSER_WIDTH = 1;
  parameter C_M_AXI_GMEM_COUT_ARUSER_WIDTH = 1;
  parameter C_M_AXI_GMEM_COUT_WUSER_WIDTH = 1;
  parameter C_M_AXI_GMEM_COUT_RUSER_WIDTH = 1;
  parameter C_M_AXI_GMEM_COUT_BUSER_WIDTH = 1;
  parameter C_M_AXI_GMEM_COUT_USER_VALUE = 0;
  parameter C_M_AXI_GMEM_COUT_PROT_VALUE = 0;
  parameter C_M_AXI_GMEM_COUT_CACHE_VALUE = 3;
  parameter C_M_AXI_GMEM_W_ID_WIDTH = 1;
  parameter C_M_AXI_GMEM_W_ADDR_WIDTH = 64;
  parameter C_M_AXI_GMEM_W_DATA_WIDTH = 512;
  parameter C_M_AXI_GMEM_W_AWUSER_WIDTH = 1;
  parameter C_M_AXI_GMEM_W_ARUSER_WIDTH = 1;
  parameter C_M_AXI_GMEM_W_WUSER_WIDTH = 1;
  parameter C_M_AXI_GMEM_W_RUSER_WIDTH = 1;
  parameter C_M_AXI_GMEM_W_BUSER_WIDTH = 1;
  parameter C_M_AXI_GMEM_W_USER_VALUE = 0;
  parameter C_M_AXI_GMEM_W_PROT_VALUE = 0;
  parameter C_M_AXI_GMEM_W_CACHE_VALUE = 3;
  parameter C_S_AXI_CONTROL_WSTRB_WIDTH = 32 / 8;
  parameter C_S_AXI_WSTRB_WIDTH = 32 / 8;
  parameter C_M_AXI_GMEM_CIN_WSTRB_WIDTH = 512 / 8;
  parameter C_M_AXI_WSTRB_WIDTH = 32 / 8;
  parameter C_M_AXI_GMEM_COUT_WSTRB_WIDTH = 512 / 8;
  parameter C_M_AXI_GMEM_W_WSTRB_WIDTH = 512 / 8;
  wire [255:0] PE_wrapper211_U0_fifo_cin_out_V_V_din_pass_0_in;
  wire [255:0] PE_wrapper211_U0_fifo_cin_out_V_V_din_pass_1_out;
  wire fifo_cin_PE_6_1_V_V_full_n_pass_0_out;
  wire fifo_cin_PE_6_1_V_V_full_n_pass_1_in;
  wire PE_wrapper211_U0_fifo_cin_out_V_V_write_pass_0_in;
  wire PE_wrapper211_U0_fifo_cin_out_V_V_write_pass_1_out;
  wire [255:0] PE_wrapper212_U0_fifo_cin_out_V_V_din_pass_0_in;
  wire [255:0] PE_wrapper212_U0_fifo_cin_out_V_V_din_pass_1_out;
  wire fifo_cin_PE_6_2_V_V_full_n_pass_0_out;
  wire fifo_cin_PE_6_2_V_V_full_n_pass_1_in;
  wire PE_wrapper212_U0_fifo_cin_out_V_V_write_pass_0_in;
  wire PE_wrapper212_U0_fifo_cin_out_V_V_write_pass_1_out;
  wire [255:0] PE_wrapper213_U0_fifo_cin_out_V_V_din_pass_0_in;
  wire [255:0] PE_wrapper213_U0_fifo_cin_out_V_V_din_pass_1_out;
  wire fifo_cin_PE_6_3_V_V_full_n_pass_0_out;
  wire fifo_cin_PE_6_3_V_V_full_n_pass_1_in;
  wire PE_wrapper213_U0_fifo_cin_out_V_V_write_pass_0_in;
  wire PE_wrapper213_U0_fifo_cin_out_V_V_write_pass_1_out;
  wire [255:0] cin_IO_L2_in125_U0_fifo_cin_out_V_V_din_pass_0_in;
  wire [255:0] cin_IO_L2_in125_U0_fifo_cin_out_V_V_din_pass_1_out;
  wire fifo_cin_cin_IO_L2_in_2_V_V_full_n_pass_0_out;
  wire fifo_cin_cin_IO_L2_in_2_V_V_full_n_pass_1_in;
  wire cin_IO_L2_in125_U0_fifo_cin_out_V_V_write_pass_0_in;
  wire cin_IO_L2_in125_U0_fifo_cin_out_V_V_write_pass_1_out;
  wire [63:0] cout_drain_IO_L1_out_wrapper424_U0_fifo_cout_drain_out_V_V_din_pass_0_in;
  wire [63:0] cout_drain_IO_L1_out_wrapper424_U0_fifo_cout_drain_out_V_V_din_pass_1_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_3_6_V_V_full_n_pass_0_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_3_6_V_V_full_n_pass_1_in;
  wire cout_drain_IO_L1_out_wrapper424_U0_fifo_cout_drain_out_V_V_write_pass_0_in;
  wire cout_drain_IO_L1_out_wrapper424_U0_fifo_cout_drain_out_V_V_write_pass_1_out;
  wire [63:0] cout_drain_IO_L1_out_wrapper408_U0_fifo_cout_drain_out_V_V_din_pass_0_in;
  wire [63:0] cout_drain_IO_L1_out_wrapper408_U0_fifo_cout_drain_out_V_V_din_pass_1_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_2_6_V_V_full_n_pass_0_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_2_6_V_V_full_n_pass_1_in;
  wire cout_drain_IO_L1_out_wrapper408_U0_fifo_cout_drain_out_V_V_write_pass_0_in;
  wire cout_drain_IO_L1_out_wrapper408_U0_fifo_cout_drain_out_V_V_write_pass_1_out;
  wire [63:0] cout_drain_IO_L1_out_wrapper376_U0_fifo_cout_drain_out_V_V_din_pass_0_in;
  wire [63:0] cout_drain_IO_L1_out_wrapper376_U0_fifo_cout_drain_out_V_V_din_pass_1_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_0_6_V_V_full_n_pass_0_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_0_6_V_V_full_n_pass_1_in;
  wire cout_drain_IO_L1_out_wrapper376_U0_fifo_cout_drain_out_V_V_write_pass_0_in;
  wire cout_drain_IO_L1_out_wrapper376_U0_fifo_cout_drain_out_V_V_write_pass_1_out;
  wire [63:0] cout_drain_IO_L1_out_wrapper392_U0_fifo_cout_drain_out_V_V_din_pass_0_in;
  wire [63:0] cout_drain_IO_L1_out_wrapper392_U0_fifo_cout_drain_out_V_V_din_pass_1_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_1_6_V_V_full_n_pass_0_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_1_6_V_V_full_n_pass_1_in;
  wire cout_drain_IO_L1_out_wrapper392_U0_fifo_cout_drain_out_V_V_write_pass_0_in;
  wire cout_drain_IO_L1_out_wrapper392_U0_fifo_cout_drain_out_V_V_write_pass_1_out;
  wire [255:0] PE_wrapper213_U0_fifo_w_out_V_V_din_pass_0_in;
  wire [255:0] PE_wrapper213_U0_fifo_w_out_V_V_din_pass_1_out;
  wire fifo_w_PE_5_4_V_V_full_n_pass_0_out;
  wire fifo_w_PE_5_4_V_V_full_n_pass_1_in;
  wire PE_wrapper213_U0_fifo_w_out_V_V_write_pass_0_in;
  wire PE_wrapper213_U0_fifo_w_out_V_V_write_pass_1_out;
  wire [255:0] PE_wrapper187_U0_fifo_w_out_V_V_din_pass_0_out;
  wire fifo_w_PE_3_2_V_V_full_n_pass_0_in;
  wire PE_wrapper187_U0_fifo_w_out_V_V_write_pass_0_out;
  wire [31:0] PE_wrapper187_U0_fifo_cout_drain_out_V_din_pass_0_out;
  wire fifo_cout_drain_PE_3_1_V_full_n_pass_0_in;
  wire PE_wrapper187_U0_fifo_cout_drain_out_V_write_pass_0_out;
  wire [255:0] PE_wrapper162_U0_fifo_cin_out_V_V_din_pass_0_in;
  wire fifo_cin_PE_2_0_V_V_full_n_pass_0_out;
  wire PE_wrapper162_U0_fifo_cin_out_V_V_write_pass_0_in;
  wire [255:0] w_IO_L2_in137_U0_fifo_w_out_V_V_din_pass_0_out;
  wire fifo_w_w_IO_L2_in_3_V_V_full_n_pass_0_in;
  wire w_IO_L2_in137_U0_fifo_w_out_V_V_write_pass_0_out;
  wire [31:0] PE_wrapper151_U0_fifo_cout_drain_out_V_din_pass_0_out;
  wire fifo_cout_drain_PE_0_1_V_full_n_pass_0_in;
  wire PE_wrapper151_U0_fifo_cout_drain_out_V_write_pass_0_out;
  wire [255:0] PE_wrapper163_U0_fifo_w_out_V_V_din_pass_0_out;
  wire fifo_w_PE_1_2_V_V_full_n_pass_0_in;
  wire PE_wrapper163_U0_fifo_w_out_V_V_write_pass_0_out;
  wire [255:0] w_IO_L2_in136_U0_fifo_w_out_V_V_din_pass_0_in;
  wire fifo_w_w_IO_L2_in_2_V_V_full_n_pass_0_out;
  wire w_IO_L2_in136_U0_fifo_w_out_V_V_write_pass_0_in;
  wire [255:0] cin_IO_L2_in124_U0_fifo_cin_out_V_V_din_pass_0_out;
  wire fifo_cin_cin_IO_L2_in_1_V_V_full_n_pass_0_in;
  wire cin_IO_L2_in124_U0_fifo_cin_out_V_V_write_pass_0_out;
  wire [255:0] w_IO_L2_in138_U0_fifo_w_local_out_V_V_din_pass_1_in;
  wire fifo_w_PE_3_0_V_V_full_n_pass_1_out;
  wire w_IO_L2_in138_U0_fifo_w_local_out_V_V_write_pass_1_in;
  wire [63:0] kernel0_entry12_U0_w_V_out_din_pass_0_out;
  wire w_V_c_full_n_pass_0_in;
  wire kernel0_entry12_U0_w_V_out_write_pass_0_out;
  wire [31:0] PE_wrapper163_U0_fifo_cout_drain_out_V_din_pass_0_out;
  wire fifo_cout_drain_PE_1_1_V_full_n_pass_0_in;
  wire PE_wrapper163_U0_fifo_cout_drain_out_V_write_pass_0_out;
  wire [255:0] PE_wrapper151_U0_fifo_w_out_V_V_din_pass_0_out;
  wire fifo_w_PE_0_2_V_V_full_n_pass_0_in;
  wire PE_wrapper151_U0_fifo_w_out_V_V_write_pass_0_out;
  wire [31:0] PE_wrapper162_U0_fifo_cout_drain_out_V_din_pass_0_in;
  wire fifo_cout_drain_PE_1_0_V_full_n_pass_0_out;
  wire PE_wrapper162_U0_fifo_cout_drain_out_V_write_pass_0_in;
  wire [255:0] PE_wrapper150_U0_fifo_cin_out_V_V_din_pass_0_out;
  wire fifo_cin_PE_1_0_V_V_full_n_pass_0_in;
  wire PE_wrapper150_U0_fifo_cin_out_V_V_write_pass_0_out;
  wire [31:0] PE_wrapper175_U0_fifo_cout_drain_out_V_din_pass_0_out;
  wire fifo_cout_drain_PE_2_1_V_full_n_pass_0_in;
  wire PE_wrapper175_U0_fifo_cout_drain_out_V_write_pass_0_out;
  wire [255:0] PE_wrapper175_U0_fifo_w_out_V_V_din_pass_0_out;
  wire fifo_w_PE_2_2_V_V_full_n_pass_0_in;
  wire PE_wrapper175_U0_fifo_w_out_V_V_write_pass_0_out;
  wire [255:0] cin_IO_L2_in125_U0_fifo_cin_local_out_V_V_din_pass_0_in;
  wire fifo_cin_PE_0_1_V_V_full_n_pass_0_out;
  wire cin_IO_L2_in125_U0_fifo_cin_local_out_V_V_write_pass_0_in;
  wire [63:0] cout_drain_IO_L1_out_wrapper378_U0_fifo_cout_drain_out_V_V_din_pass_1_in;
  wire fifo_cout_drain_cout_drain_IO_L1_out_0_4_V_V_full_n_pass_1_out;
  wire cout_drain_IO_L1_out_wrapper378_U0_fifo_cout_drain_out_V_V_write_pass_1_in;
  wire [63:0] kernel0_entry12_U0_cout_V_out_din_pass_0_out;
  wire cout_V_c_full_n_pass_0_in;
  wire kernel0_entry12_U0_cout_V_out_write_pass_0_out;
  wire [255:0] PE_wrapper187_U0_fifo_cin_out_V_V_din_pass_0_out;
  wire fifo_cin_PE_4_1_V_V_full_n_pass_0_in;
  wire PE_wrapper187_U0_fifo_cin_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper162_U0_fifo_w_out_V_V_din_pass_0_in;
  wire fifo_w_PE_1_1_V_V_full_n_pass_0_out;
  wire PE_wrapper162_U0_fifo_w_out_V_V_write_pass_0_in;
  wire [63:0] cout_drain_IO_L1_out_wrapper382_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_0_0_V_V_full_n_pass_0_in;
  wire cout_drain_IO_L1_out_wrapper382_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper186_U0_fifo_cin_out_V_V_din_pass_0_out;
  wire fifo_cin_PE_4_0_V_V_full_n_pass_0_in;
  wire PE_wrapper186_U0_fifo_cin_out_V_V_write_pass_0_out;
  wire [255:0] w_IO_L2_in135_U0_fifo_w_local_out_V_V_din_pass_0_in;
  wire fifo_w_PE_0_0_V_V_full_n_pass_0_out;
  wire w_IO_L2_in135_U0_fifo_w_local_out_V_V_write_pass_0_in;
  wire ap_start_Boundary_X4Y2_To_X6Y2_out;
  wire ap_rst_n_Boundary_X4Y2_To_X6Y2_out;
  wire ap_done_Boundary_X4Y2_To_X6Y2_in;
  wire ap_start_Boundary_X6Y0_To_X6Y2_out;
  wire ap_rst_n_Boundary_X6Y0_To_X6Y2_out;
  wire ap_done_Boundary_X6Y0_To_X6Y2_in;
  wire ap_start_Boundary_X4Y0_To_X4Y2_out;
  wire ap_rst_n_Boundary_X4Y0_To_X4Y2_out;
  wire ap_done_Boundary_X4Y0_To_X4Y2_in;
  wire [255:0] PE_wrapper190_U0_fifo_w_out_V_V_din_pass_0_in;
  wire [255:0] PE_wrapper190_U0_fifo_w_out_V_V_din_pass_1_out;
  wire fifo_w_PE_3_5_V_V_full_n_pass_0_out;
  wire fifo_w_PE_3_5_V_V_full_n_pass_1_in;
  wire PE_wrapper190_U0_fifo_w_out_V_V_write_pass_0_in;
  wire PE_wrapper190_U0_fifo_w_out_V_V_write_pass_1_out;
  wire [255:0] PE_wrapper179_U0_fifo_cin_out_V_V_din_pass_0_in;
  wire [255:0] PE_wrapper179_U0_fifo_cin_out_V_V_din_pass_1_out;
  wire fifo_cin_PE_3_5_V_V_full_n_pass_0_out;
  wire fifo_cin_PE_3_5_V_V_full_n_pass_1_in;
  wire PE_wrapper179_U0_fifo_cin_out_V_V_write_pass_0_in;
  wire PE_wrapper179_U0_fifo_cin_out_V_V_write_pass_1_out;
  wire [63:0] kernel0_entry12_U0_cout_V_out_din_pass_1_in;
  wire [63:0] kernel0_entry12_U0_cout_V_out_din_pass_2_out;
  wire cout_V_c_full_n_pass_1_out;
  wire cout_V_c_full_n_pass_2_in;
  wire kernel0_entry12_U0_cout_V_out_write_pass_1_in;
  wire kernel0_entry12_U0_cout_V_out_write_pass_2_out;
  wire [255:0] PE_wrapper190_U0_fifo_cin_out_V_V_din_pass_0_in;
  wire fifo_cin_PE_4_4_V_V_full_n_pass_0_out;
  wire PE_wrapper190_U0_fifo_cin_out_V_V_write_pass_0_in;
  wire [255:0] PE_wrapper201_U0_fifo_w_out_V_V_din_pass_1_in;
  wire fifo_w_PE_4_4_V_V_full_n_pass_1_out;
  wire PE_wrapper201_U0_fifo_w_out_V_V_write_pass_1_in;
  wire [63:0] cout_drain_IO_L1_out_wrapper440_U0_fifo_cout_drain_out_V_V_din_pass_1_in;
  wire fifo_cout_drain_cout_drain_IO_L1_out_4_6_V_V_full_n_pass_1_out;
  wire cout_drain_IO_L1_out_wrapper440_U0_fifo_cout_drain_out_V_V_write_pass_1_in;
  wire [255:0] PE_wrapper213_U0_fifo_w_out_V_V_din_pass_2_in;
  wire fifo_w_PE_5_4_V_V_full_n_pass_2_out;
  wire PE_wrapper213_U0_fifo_w_out_V_V_write_pass_2_in;
  wire [255:0] PE_wrapper214_U0_fifo_w_out_V_V_din_pass_0_out;
  wire fifo_w_PE_5_5_V_V_full_n_pass_0_in;
  wire PE_wrapper214_U0_fifo_w_out_V_V_write_pass_0_out;
  wire [63:0] cout_drain_IO_L1_out_wrapper441_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_4_5_V_V_full_n_pass_0_in;
  wire cout_drain_IO_L1_out_wrapper441_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  wire [255:0] w_IO_L3_in_serialize_U0_fifo_w_local_out_V_V_din_pass_0_out;
  wire fifo_w_w_IO_L3_in_serialize_V_V_full_n_pass_0_in;
  wire w_IO_L3_in_serialize_U0_fifo_w_local_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper214_U0_fifo_cin_out_V_V_din_pass_0_out;
  wire fifo_cin_PE_6_4_V_V_full_n_pass_0_in;
  wire PE_wrapper214_U0_fifo_cin_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper202_U0_fifo_w_out_V_V_din_pass_0_out;
  wire fifo_w_PE_4_5_V_V_full_n_pass_0_in;
  wire PE_wrapper202_U0_fifo_w_out_V_V_write_pass_0_out;
  wire [31:0] PE_wrapper202_U0_fifo_cout_drain_out_V_din_pass_0_out;
  wire fifo_cout_drain_PE_4_4_V_full_n_pass_0_in;
  wire PE_wrapper202_U0_fifo_cout_drain_out_V_write_pass_0_out;
  wire [63:0] kernel0_entry12_U0_w_V_out_din_pass_1_in;
  wire w_V_c_full_n_pass_1_out;
  wire kernel0_entry12_U0_w_V_out_write_pass_1_in;
  wire ap_start_Boundary_X4Y4_To_X6Y4_in;
  wire ap_rst_n_Boundary_X4Y4_To_X6Y4_in;
  wire ap_done_Boundary_X4Y4_To_X6Y4_out;
  wire ap_start_Boundary_X4Y6_To_X6Y6_out;
  wire ap_rst_n_Boundary_X4Y6_To_X6Y6_out;
  wire ap_done_Boundary_X4Y6_To_X6Y6_in;
  wire [255:0] PE_wrapper230_U0_fifo_w_out_V_V_din_pass_0_in;
  wire [255:0] PE_wrapper230_U0_fifo_w_out_V_V_din_pass_1_out;
  wire fifo_w_PE_6_9_V_V_full_n_pass_0_out;
  wire fifo_w_PE_6_9_V_V_full_n_pass_1_in;
  wire PE_wrapper230_U0_fifo_w_out_V_V_write_pass_0_in;
  wire PE_wrapper230_U0_fifo_w_out_V_V_write_pass_1_out;
  wire [63:0] cout_drain_IO_L1_out_wrapper522_U0_fifo_cout_drain_out_V_V_din_pass_0_in;
  wire [63:0] cout_drain_IO_L1_out_wrapper522_U0_fifo_cout_drain_out_V_V_din_pass_1_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_9_4_V_V_full_n_pass_0_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_9_4_V_V_full_n_pass_1_in;
  wire cout_drain_IO_L1_out_wrapper522_U0_fifo_cout_drain_out_V_V_write_pass_0_in;
  wire cout_drain_IO_L1_out_wrapper522_U0_fifo_cout_drain_out_V_V_write_pass_1_out;
  wire [63:0] cout_drain_IO_L1_out_wrapper542_U0_fifo_cout_drain_out_V_V_din_pass_0_in;
  wire [63:0] cout_drain_IO_L1_out_wrapper542_U0_fifo_cout_drain_out_V_V_din_pass_1_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_10_0_V_V_full_n_pass_0_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_10_0_V_V_full_n_pass_1_in;
  wire cout_drain_IO_L1_out_wrapper542_U0_fifo_cout_drain_out_V_V_write_pass_0_in;
  wire cout_drain_IO_L1_out_wrapper542_U0_fifo_cout_drain_out_V_V_write_pass_1_out;
  wire [255:0] PE_wrapper219_U0_fifo_cin_out_V_V_din_pass_0_in;
  wire [255:0] PE_wrapper219_U0_fifo_cin_out_V_V_din_pass_1_out;
  wire fifo_cin_PE_6_9_V_V_full_n_pass_0_out;
  wire fifo_cin_PE_6_9_V_V_full_n_pass_1_in;
  wire PE_wrapper219_U0_fifo_cin_out_V_V_write_pass_0_in;
  wire PE_wrapper219_U0_fifo_cin_out_V_V_write_pass_1_out;
  wire [255:0] PE_wrapper172_U0_fifo_cin_out_V_V_din_pass_0_in;
  wire [255:0] PE_wrapper172_U0_fifo_cin_out_V_V_din_pass_1_out;
  wire fifo_cin_PE_2_10_V_V_full_n_pass_0_out;
  wire fifo_cin_PE_2_10_V_V_full_n_pass_1_in;
  wire PE_wrapper172_U0_fifo_cin_out_V_V_write_pass_0_in;
  wire PE_wrapper172_U0_fifo_cin_out_V_V_write_pass_1_out;
  wire [255:0] cin_IO_L2_in134_U0_fifo_cin_out_V_V_din_pass_0_in;
  wire [255:0] cin_IO_L2_in134_U0_fifo_cin_out_V_V_din_pass_1_out;
  wire fifo_cin_cin_IO_L2_in_11_V_V_full_n_pass_0_out;
  wire fifo_cin_cin_IO_L2_in_11_V_V_full_n_pass_1_in;
  wire cin_IO_L2_in134_U0_fifo_cin_out_V_V_write_pass_0_in;
  wire cin_IO_L2_in134_U0_fifo_cin_out_V_V_write_pass_1_out;
  wire [255:0] PE_wrapper194_U0_fifo_w_out_V_V_din_pass_1_in;
  wire [255:0] PE_wrapper194_U0_fifo_w_out_V_V_din_pass_2_out;
  wire fifo_w_PE_3_9_V_V_full_n_pass_1_out;
  wire fifo_w_PE_3_9_V_V_full_n_pass_2_in;
  wire PE_wrapper194_U0_fifo_w_out_V_V_write_pass_1_in;
  wire PE_wrapper194_U0_fifo_w_out_V_V_write_pass_2_out;
  wire [63:0] cout_drain_IO_L1_out_wrapper548_U0_fifo_cout_drain_out_V_V_din_pass_0_in;
  wire [63:0] cout_drain_IO_L1_out_wrapper548_U0_fifo_cout_drain_out_V_V_din_pass_1_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_11_9_V_V_full_n_pass_0_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_11_9_V_V_full_n_pass_1_in;
  wire cout_drain_IO_L1_out_wrapper548_U0_fifo_cout_drain_out_V_V_write_pass_0_in;
  wire cout_drain_IO_L1_out_wrapper548_U0_fifo_cout_drain_out_V_V_write_pass_1_out;
  wire [31:0] PE_wrapper219_U0_fifo_cout_drain_out_V_din_pass_0_in;
  wire [31:0] PE_wrapper219_U0_fifo_cout_drain_out_V_din_pass_1_out;
  wire fifo_cout_drain_PE_5_9_V_full_n_pass_0_out;
  wire fifo_cout_drain_PE_5_9_V_full_n_pass_1_in;
  wire PE_wrapper219_U0_fifo_cout_drain_out_V_write_pass_0_in;
  wire PE_wrapper219_U0_fifo_cout_drain_out_V_write_pass_1_out;
  wire [63:0] cout_drain_IO_L1_out_wrapper517_U0_fifo_cout_drain_out_V_V_din_pass_0_in;
  wire [63:0] cout_drain_IO_L1_out_wrapper517_U0_fifo_cout_drain_out_V_V_din_pass_1_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_9_9_V_V_full_n_pass_0_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_9_9_V_V_full_n_pass_1_in;
  wire cout_drain_IO_L1_out_wrapper517_U0_fifo_cout_drain_out_V_V_write_pass_0_in;
  wire cout_drain_IO_L1_out_wrapper517_U0_fifo_cout_drain_out_V_V_write_pass_1_out;
  wire [63:0] cout_drain_IO_L1_out_wrapper533_U0_fifo_cout_drain_out_V_V_din_pass_0_in;
  wire [63:0] cout_drain_IO_L1_out_wrapper533_U0_fifo_cout_drain_out_V_V_din_pass_1_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_10_9_V_V_full_n_pass_0_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_10_9_V_V_full_n_pass_1_in;
  wire cout_drain_IO_L1_out_wrapper533_U0_fifo_cout_drain_out_V_V_write_pass_0_in;
  wire cout_drain_IO_L1_out_wrapper533_U0_fifo_cout_drain_out_V_V_write_pass_1_out;
  wire [63:0] cout_drain_IO_L1_out_wrapper535_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_10_7_V_V_full_n_pass_0_in;
  wire cout_drain_IO_L1_out_wrapper535_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper219_U0_fifo_w_out_V_V_din_pass_0_in;
  wire fifo_w_PE_5_10_V_V_full_n_pass_0_out;
  wire PE_wrapper219_U0_fifo_w_out_V_V_write_pass_0_in;
  wire [63:0] cout_drain_IO_L1_out_wrapper537_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_10_5_V_V_full_n_pass_0_in;
  wire cout_drain_IO_L1_out_wrapper537_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper171_U0_fifo_cin_out_V_V_din_pass_0_in;
  wire fifo_cin_PE_2_9_V_V_full_n_pass_0_out;
  wire PE_wrapper171_U0_fifo_cin_out_V_V_write_pass_0_in;
  wire [255:0] PE_wrapper172_U0_fifo_w_out_V_V_din_pass_0_in;
  wire fifo_w_PE_1_11_V_V_full_n_pass_0_out;
  wire PE_wrapper172_U0_fifo_w_out_V_V_write_pass_0_in;
  wire [63:0] cout_drain_IO_L1_out_wrapper551_U0_fifo_cout_drain_out_V_V_din_pass_1_in;
  wire fifo_cout_drain_cout_drain_IO_L1_out_11_6_V_V_full_n_pass_1_out;
  wire cout_drain_IO_L1_out_wrapper551_U0_fifo_cout_drain_out_V_V_write_pass_1_in;
  wire [63:0] cout_drain_IO_L1_out_wrapper555_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_11_2_V_V_full_n_pass_0_in;
  wire cout_drain_IO_L1_out_wrapper555_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper196_U0_fifo_cin_out_V_V_din_pass_0_in;
  wire fifo_cin_PE_4_10_V_V_full_n_pass_0_out;
  wire PE_wrapper196_U0_fifo_cin_out_V_V_write_pass_0_in;
  wire [63:0] cout_drain_IO_L1_out_wrapper539_U0_fifo_cout_drain_out_V_V_din_pass_0_in;
  wire fifo_cout_drain_cout_drain_IO_L1_out_10_3_V_V_full_n_pass_0_out;
  wire cout_drain_IO_L1_out_wrapper539_U0_fifo_cout_drain_out_V_V_write_pass_0_in;
  wire [255:0] PE_wrapper244_U0_fifo_cin_out_V_V_din_pass_0_out;
  wire fifo_cin_PE_8_10_V_V_full_n_pass_0_in;
  wire PE_wrapper244_U0_fifo_cin_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper231_U0_fifo_w_out_V_V_din_pass_0_in;
  wire fifo_w_PE_6_10_V_V_full_n_pass_0_out;
  wire PE_wrapper231_U0_fifo_w_out_V_V_write_pass_0_in;
  wire [255:0] PE_wrapper173_U0_fifo_w_out_V_V_din_pass_0_out;
  wire fifo_w_PE_1_12_V_V_full_n_pass_0_in;
  wire PE_wrapper173_U0_fifo_w_out_V_V_write_pass_0_out;
  wire [31:0] PE_wrapper231_U0_fifo_cout_drain_out_V_din_pass_0_in;
  wire fifo_cout_drain_PE_6_9_V_full_n_pass_0_out;
  wire PE_wrapper231_U0_fifo_cout_drain_out_V_write_pass_0_in;
  wire [255:0] PE_wrapper207_U0_fifo_w_out_V_V_din_pass_0_in;
  wire fifo_w_PE_4_10_V_V_full_n_pass_0_out;
  wire PE_wrapper207_U0_fifo_w_out_V_V_write_pass_0_in;
  wire [31:0] PE_wrapper221_U0_fifo_cout_drain_out_V_din_pass_0_in;
  wire fifo_cout_drain_PE_5_11_V_full_n_pass_0_out;
  wire PE_wrapper221_U0_fifo_cout_drain_out_V_write_pass_0_in;
  wire [31:0] PE_wrapper183_U0_fifo_cout_drain_out_V_din_pass_0_out;
  wire fifo_cout_drain_PE_2_9_V_full_n_pass_0_in;
  wire PE_wrapper183_U0_fifo_cout_drain_out_V_write_pass_0_out;
  wire [255:0] PE_wrapper161_U0_fifo_cin_out_V_V_din_pass_1_in;
  wire fifo_cin_PE_1_11_V_V_full_n_pass_1_out;
  wire PE_wrapper161_U0_fifo_cin_out_V_V_write_pass_1_in;
  wire [31:0] PE_wrapper232_U0_fifo_cout_drain_out_V_din_pass_0_out;
  wire fifo_cout_drain_PE_6_10_V_full_n_pass_0_in;
  wire PE_wrapper232_U0_fifo_cout_drain_out_V_write_pass_0_out;
  wire [63:0] kernel0_entry12_U0_cout_V_out_din_pass_5_in;
  wire cout_V_c_full_n_pass_5_out;
  wire kernel0_entry12_U0_cout_V_out_write_pass_5_in;
  wire [63:0] cout_drain_IO_L1_out_wrapper540_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_10_2_V_V_full_n_pass_0_in;
  wire cout_drain_IO_L1_out_wrapper540_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  wire [63:0] cout_drain_IO_L1_out_wrapper552_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_11_5_V_V_full_n_pass_0_in;
  wire cout_drain_IO_L1_out_wrapper552_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper243_U0_fifo_w_out_V_V_din_pass_3_in;
  wire fifo_w_PE_7_10_V_V_full_n_pass_3_out;
  wire PE_wrapper243_U0_fifo_w_out_V_V_write_pass_3_in;
  wire [31:0] PE_wrapper243_U0_fifo_cout_drain_out_V_din_pass_3_in;
  wire fifo_cout_drain_PE_7_9_V_full_n_pass_3_out;
  wire PE_wrapper243_U0_fifo_cout_drain_out_V_write_pass_3_in;
  wire [31:0] PE_wrapper184_U0_fifo_cout_drain_out_V_din_pass_0_in;
  wire fifo_cout_drain_PE_2_10_V_full_n_pass_0_out;
  wire PE_wrapper184_U0_fifo_cout_drain_out_V_write_pass_0_in;
  wire [255:0] PE_wrapper243_U0_fifo_cin_out_V_V_din_pass_3_in;
  wire fifo_cin_PE_8_9_V_V_full_n_pass_3_out;
  wire PE_wrapper243_U0_fifo_cin_out_V_V_write_pass_3_in;
  wire [31:0] PE_wrapper255_U0_fifo_cout_drain_out_V_din_pass_0_out;
  wire fifo_cout_drain_PE_8_9_V_full_n_pass_0_in;
  wire PE_wrapper255_U0_fifo_cout_drain_out_V_write_pass_0_out;
  wire [31:0] PE_wrapper185_U0_fifo_cout_drain_out_V_din_pass_1_in;
  wire fifo_cout_drain_PE_2_11_V_full_n_pass_1_out;
  wire PE_wrapper185_U0_fifo_cout_drain_out_V_write_pass_1_in;
  wire [63:0] cout_drain_IO_L1_out_wrapper518_U0_fifo_cout_drain_out_V_V_din_pass_1_in;
  wire fifo_cout_drain_cout_drain_IO_L1_out_9_8_V_V_full_n_pass_1_out;
  wire cout_drain_IO_L1_out_wrapper518_U0_fifo_cout_drain_out_V_V_write_pass_1_in;
  wire [255:0] PE_wrapper255_U0_fifo_cin_out_V_V_din_pass_0_out;
  wire fifo_cin_PE_9_9_V_V_full_n_pass_0_in;
  wire PE_wrapper255_U0_fifo_cin_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper244_U0_fifo_w_out_V_V_din_pass_0_out;
  wire fifo_w_PE_7_11_V_V_full_n_pass_0_in;
  wire PE_wrapper244_U0_fifo_w_out_V_V_write_pass_0_out;
  wire [31:0] PE_wrapper173_U0_fifo_cout_drain_out_V_din_pass_0_out;
  wire fifo_cout_drain_PE_1_11_V_full_n_pass_0_in;
  wire PE_wrapper173_U0_fifo_cout_drain_out_V_write_pass_0_out;
  wire [255:0] PE_wrapper254_U0_fifo_w_out_V_V_din_pass_0_in;
  wire fifo_w_PE_8_9_V_V_full_n_pass_0_out;
  wire PE_wrapper254_U0_fifo_w_out_V_V_write_pass_0_in;
  wire [31:0] PE_wrapper208_U0_fifo_cout_drain_out_V_din_pass_0_out;
  wire fifo_cout_drain_PE_4_10_V_full_n_pass_0_in;
  wire PE_wrapper208_U0_fifo_cout_drain_out_V_write_pass_0_out;
  wire [63:0] cout_drain_IO_L1_out_wrapper536_U0_fifo_cout_drain_out_V_V_din_pass_0_in;
  wire fifo_cout_drain_cout_drain_IO_L1_out_10_6_V_V_full_n_pass_0_out;
  wire cout_drain_IO_L1_out_wrapper536_U0_fifo_cout_drain_out_V_V_write_pass_0_in;
  wire [255:0] PE_wrapper182_U0_fifo_w_out_V_V_din_pass_1_in;
  wire fifo_w_PE_2_9_V_V_full_n_pass_1_out;
  wire PE_wrapper182_U0_fifo_w_out_V_V_write_pass_1_in;
  wire [255:0] PE_wrapper220_U0_fifo_w_out_V_V_din_pass_0_out;
  wire fifo_w_PE_5_11_V_V_full_n_pass_0_in;
  wire PE_wrapper220_U0_fifo_w_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper255_U0_fifo_w_out_V_V_din_pass_0_out;
  wire fifo_w_PE_8_10_V_V_full_n_pass_0_in;
  wire PE_wrapper255_U0_fifo_w_out_V_V_write_pass_0_out;
  wire [63:0] cout_drain_IO_L1_out_wrapper534_U0_fifo_cout_drain_out_V_V_din_pass_1_in;
  wire fifo_cout_drain_cout_drain_IO_L1_out_10_8_V_V_full_n_pass_1_out;
  wire cout_drain_IO_L1_out_wrapper534_U0_fifo_cout_drain_out_V_V_write_pass_1_in;
  wire [63:0] cout_drain_IO_L1_out_wrapper520_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_9_6_V_V_full_n_pass_0_in;
  wire cout_drain_IO_L1_out_wrapper520_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  wire [63:0] cout_drain_IO_L3_out_U0_fifo_cout_drain_out_V_V_din_pass_2_in;
  wire fifo_cout_drain_cout_drain_IO_L3_out_serialize_V_V_full_n_pass_2_out;
  wire cout_drain_IO_L3_out_U0_fifo_cout_drain_out_V_V_write_pass_2_in;
  wire [255:0] PE_wrapper173_U0_fifo_cin_out_V_V_din_pass_0_out;
  wire fifo_cin_PE_2_11_V_V_full_n_pass_0_in;
  wire PE_wrapper173_U0_fifo_cin_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper232_U0_fifo_w_out_V_V_din_pass_0_out;
  wire fifo_w_PE_6_11_V_V_full_n_pass_0_in;
  wire PE_wrapper232_U0_fifo_w_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper183_U0_fifo_w_out_V_V_din_pass_0_out;
  wire fifo_w_PE_2_10_V_V_full_n_pass_0_in;
  wire PE_wrapper183_U0_fifo_w_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper221_U0_fifo_w_out_V_V_din_pass_0_in;
  wire fifo_w_PE_5_12_V_V_full_n_pass_0_out;
  wire PE_wrapper221_U0_fifo_w_out_V_V_write_pass_0_in;
  wire [255:0] PE_wrapper208_U0_fifo_w_out_V_V_din_pass_0_out;
  wire fifo_w_PE_4_11_V_V_full_n_pass_0_in;
  wire PE_wrapper208_U0_fifo_w_out_V_V_write_pass_0_out;
  wire [31:0] PE_wrapper197_U0_fifo_cout_drain_out_V_din_pass_1_in;
  wire fifo_cout_drain_PE_3_11_V_full_n_pass_1_out;
  wire PE_wrapper197_U0_fifo_cout_drain_out_V_write_pass_1_in;
  wire [255:0] PE_wrapper183_U0_fifo_cin_out_V_V_din_pass_0_out;
  wire fifo_cin_PE_3_9_V_V_full_n_pass_0_in;
  wire PE_wrapper183_U0_fifo_cin_out_V_V_write_pass_0_out;
  wire [63:0] cout_drain_IO_L1_out_wrapper553_U0_fifo_cout_drain_out_V_V_din_pass_0_in;
  wire fifo_cout_drain_cout_drain_IO_L1_out_11_4_V_V_full_n_pass_0_out;
  wire cout_drain_IO_L1_out_wrapper553_U0_fifo_cout_drain_out_V_V_write_pass_0_in;
  wire ap_start_Boundary_X4Y12_To_X6Y12_in;
  wire ap_rst_n_Boundary_X4Y12_To_X6Y12_in;
  wire ap_done_Boundary_X4Y12_To_X6Y12_out;
  wire ap_start_Boundary_X4Y14_To_X6Y14_out;
  wire ap_rst_n_Boundary_X4Y14_To_X6Y14_out;
  wire ap_done_Boundary_X4Y14_To_X6Y14_in;
  wire [255:0] PE_wrapper260_U0_fifo_cin_out_V_V_din_pass_0_in;
  wire [255:0] PE_wrapper260_U0_fifo_cin_out_V_V_din_pass_1_out;
  wire fifo_cin_PE_10_2_V_V_full_n_pass_0_out;
  wire fifo_cin_PE_10_2_V_V_full_n_pass_1_in;
  wire PE_wrapper260_U0_fifo_cin_out_V_V_write_pass_0_in;
  wire PE_wrapper260_U0_fifo_cin_out_V_V_write_pass_1_out;
  wire [255:0] PE_wrapper261_U0_fifo_w_out_V_V_din_pass_0_in;
  wire [255:0] PE_wrapper261_U0_fifo_w_out_V_V_din_pass_1_out;
  wire fifo_w_PE_9_4_V_V_full_n_pass_0_out;
  wire fifo_w_PE_9_4_V_V_full_n_pass_1_in;
  wire PE_wrapper261_U0_fifo_w_out_V_V_write_pass_0_in;
  wire PE_wrapper261_U0_fifo_w_out_V_V_write_pass_1_out;
  wire [255:0] w_IO_L2_in144_U0_fifo_w_out_V_V_din_pass_0_out;
  wire fifo_w_w_IO_L2_in_10_V_V_full_n_pass_0_in;
  wire w_IO_L2_in144_U0_fifo_w_out_V_V_write_pass_0_out;
  wire [31:0] PE_wrapper271_U0_fifo_cout_drain_out_V_din_pass_0_out;
  wire fifo_cout_drain_PE_10_1_V_full_n_pass_0_in;
  wire PE_wrapper271_U0_fifo_cout_drain_out_V_write_pass_0_out;
  wire [63:0] cout_drain_IO_L1_out_wrapper372_U0_fifo_cout_drain_out_V_V_din_pass_0_in;
  wire fifo_cout_drain_cout_drain_IO_L1_out_0_10_V_V_full_n_pass_0_out;
  wire cout_drain_IO_L1_out_wrapper372_U0_fifo_cout_drain_out_V_V_write_pass_0_in;
  wire [31:0] PE_wrapper247_U0_fifo_cout_drain_out_V_din_pass_0_out;
  wire fifo_cout_drain_PE_8_1_V_full_n_pass_0_in;
  wire PE_wrapper247_U0_fifo_cout_drain_out_V_write_pass_0_out;
  wire [31:0] PE_wrapper259_U0_fifo_cout_drain_out_V_din_pass_0_out;
  wire fifo_cout_drain_PE_9_1_V_full_n_pass_0_in;
  wire PE_wrapper259_U0_fifo_cout_drain_out_V_write_pass_0_out;
  wire [255:0] PE_wrapper234_U0_fifo_cin_out_V_V_din_pass_1_in;
  wire fifo_cin_PE_8_0_V_V_full_n_pass_1_out;
  wire PE_wrapper234_U0_fifo_cin_out_V_V_write_pass_1_in;
  wire [255:0] PE_wrapper258_U0_fifo_cin_out_V_V_din_pass_0_out;
  wire fifo_cin_PE_10_0_V_V_full_n_pass_0_in;
  wire PE_wrapper258_U0_fifo_cin_out_V_V_write_pass_0_out;
  wire [63:0] cout_drain_IO_L1_out_wrapper374_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_0_8_V_V_full_n_pass_0_in;
  wire cout_drain_IO_L1_out_wrapper374_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper235_U0_fifo_cin_out_V_V_din_pass_1_in;
  wire fifo_cin_PE_8_1_V_V_full_n_pass_1_out;
  wire PE_wrapper235_U0_fifo_cin_out_V_V_write_pass_1_in;
  wire [255:0] PE_wrapper247_U0_fifo_w_out_V_V_din_pass_0_out;
  wire fifo_w_PE_8_2_V_V_full_n_pass_0_in;
  wire PE_wrapper247_U0_fifo_w_out_V_V_write_pass_0_out;
  wire [255:0] w_IO_L2_in142_U0_fifo_w_out_V_V_din_pass_1_in;
  wire fifo_w_w_IO_L2_in_8_V_V_full_n_pass_1_out;
  wire w_IO_L2_in142_U0_fifo_w_out_V_V_write_pass_1_in;
  wire [255:0] PE_wrapper271_U0_fifo_cin_out_V_V_din_pass_0_out;
  wire fifo_cin_PE_11_1_V_V_full_n_pass_0_in;
  wire PE_wrapper271_U0_fifo_cin_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper270_U0_fifo_w_out_V_V_din_pass_0_in;
  wire fifo_w_PE_10_1_V_V_full_n_pass_0_out;
  wire PE_wrapper270_U0_fifo_w_out_V_V_write_pass_0_in;
  wire [255:0] PE_wrapper259_U0_fifo_w_out_V_V_din_pass_0_out;
  wire fifo_w_PE_9_2_V_V_full_n_pass_0_in;
  wire PE_wrapper259_U0_fifo_w_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper271_U0_fifo_w_out_V_V_din_pass_0_out;
  wire fifo_w_PE_10_2_V_V_full_n_pass_0_in;
  wire PE_wrapper271_U0_fifo_w_out_V_V_write_pass_0_out;
  wire ap_start_Boundary_X2Y0_To_X2Y2_in;
  wire ap_rst_n_Boundary_X2Y0_To_X2Y2_in;
  wire ap_done_Boundary_X2Y0_To_X2Y2_out;
  wire ap_start_Boundary_X0Y2_To_X2Y2_out;
  wire ap_rst_n_Boundary_X0Y2_To_X2Y2_out;
  wire ap_done_Boundary_X0Y2_To_X2Y2_in;
  wire [255:0] PE_wrapper234_U0_fifo_cin_out_V_V_din_pass_0_in;
  wire [255:0] PE_wrapper234_U0_fifo_cin_out_V_V_din_pass_1_out;
  wire fifo_cin_PE_8_0_V_V_full_n_pass_0_out;
  wire fifo_cin_PE_8_0_V_V_full_n_pass_1_in;
  wire PE_wrapper234_U0_fifo_cin_out_V_V_write_pass_0_in;
  wire PE_wrapper234_U0_fifo_cin_out_V_V_write_pass_1_out;
  wire [255:0] PE_wrapper235_U0_fifo_cin_out_V_V_din_pass_0_in;
  wire [255:0] PE_wrapper235_U0_fifo_cin_out_V_V_din_pass_1_out;
  wire fifo_cin_PE_8_1_V_V_full_n_pass_0_out;
  wire fifo_cin_PE_8_1_V_V_full_n_pass_1_in;
  wire PE_wrapper235_U0_fifo_cin_out_V_V_write_pass_0_in;
  wire PE_wrapper235_U0_fifo_cin_out_V_V_write_pass_1_out;
  wire [255:0] w_IO_L2_in142_U0_fifo_w_out_V_V_din_pass_0_in;
  wire [255:0] w_IO_L2_in142_U0_fifo_w_out_V_V_din_pass_1_out;
  wire fifo_w_w_IO_L2_in_8_V_V_full_n_pass_0_out;
  wire fifo_w_w_IO_L2_in_8_V_V_full_n_pass_1_in;
  wire w_IO_L2_in142_U0_fifo_w_out_V_V_write_pass_0_in;
  wire w_IO_L2_in142_U0_fifo_w_out_V_V_write_pass_1_out;
  wire [255:0] PE_wrapper261_U0_fifo_w_out_V_V_din_pass_1_in;
  wire [255:0] PE_wrapper261_U0_fifo_w_out_V_V_din_pass_2_out;
  wire fifo_w_PE_9_4_V_V_full_n_pass_1_out;
  wire fifo_w_PE_9_4_V_V_full_n_pass_2_in;
  wire PE_wrapper261_U0_fifo_w_out_V_V_write_pass_1_in;
  wire PE_wrapper261_U0_fifo_w_out_V_V_write_pass_2_out;
  wire [255:0] PE_wrapper237_U0_fifo_w_out_V_V_din_pass_0_in;
  wire [255:0] PE_wrapper237_U0_fifo_w_out_V_V_din_pass_1_out;
  wire fifo_w_PE_7_4_V_V_full_n_pass_0_out;
  wire fifo_w_PE_7_4_V_V_full_n_pass_1_in;
  wire PE_wrapper237_U0_fifo_w_out_V_V_write_pass_0_in;
  wire PE_wrapper237_U0_fifo_w_out_V_V_write_pass_1_out;
  wire [255:0] PE_wrapper260_U0_fifo_cin_out_V_V_din_pass_1_in;
  wire fifo_cin_PE_10_2_V_V_full_n_pass_1_out;
  wire PE_wrapper260_U0_fifo_cin_out_V_V_write_pass_1_in;
  wire [63:0] cout_drain_IO_L1_out_wrapper402_U0_fifo_cout_drain_out_V_V_din_pass_2_in;
  wire fifo_cout_drain_cout_drain_IO_L1_out_2_12_V_V_full_n_pass_2_out;
  wire cout_drain_IO_L1_out_wrapper402_U0_fifo_cout_drain_out_V_V_write_pass_2_in;
  wire [255:0] PE_wrapper271_U0_fifo_w_out_V_V_din_pass_0_in;
  wire fifo_w_PE_10_2_V_V_full_n_pass_0_out;
  wire PE_wrapper271_U0_fifo_w_out_V_V_write_pass_0_in;
  wire [63:0] cout_drain_IO_L1_out_wrapper372_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_0_10_V_V_full_n_pass_0_in;
  wire cout_drain_IO_L1_out_wrapper372_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  wire [31:0] PE_wrapper247_U0_fifo_cout_drain_out_V_din_pass_0_in;
  wire fifo_cout_drain_PE_8_1_V_full_n_pass_0_out;
  wire PE_wrapper247_U0_fifo_cout_drain_out_V_write_pass_0_in;
  wire [255:0] PE_wrapper282_U0_fifo_cin_out_V_V_din_pass_0_out;
  wire fifo_cin_PE_12_0_V_V_full_n_pass_0_in;
  wire PE_wrapper282_U0_fifo_cin_out_V_V_write_pass_0_out;
  wire [255:0] w_IO_L2_in146_U0_fifo_w_out_V_V_din_pass_0_out;
  wire fifo_w_w_IO_L2_in_12_V_V_full_n_pass_0_in;
  wire w_IO_L2_in146_U0_fifo_w_out_V_V_write_pass_0_out;
  wire [31:0] PE_wrapper294_U0_fifo_cout_drain_out_V_din_pass_1_in;
  wire fifo_cout_drain_PE_12_0_V_full_n_pass_1_out;
  wire PE_wrapper294_U0_fifo_cout_drain_out_V_write_pass_1_in;
  wire [255:0] PE_wrapper271_U0_fifo_cin_out_V_V_din_pass_0_in;
  wire fifo_cin_PE_11_1_V_V_full_n_pass_0_out;
  wire PE_wrapper271_U0_fifo_cin_out_V_V_write_pass_0_in;
  wire [255:0] w_IO_L2_in144_U0_fifo_w_out_V_V_din_pass_0_in;
  wire fifo_w_w_IO_L2_in_10_V_V_full_n_pass_0_out;
  wire w_IO_L2_in144_U0_fifo_w_out_V_V_write_pass_0_in;
  wire [63:0] cout_drain_IO_L1_out_wrapper386_U0_fifo_cout_drain_out_V_V_din_pass_0_in;
  wire fifo_cout_drain_cout_drain_IO_L1_out_1_12_V_V_full_n_pass_0_out;
  wire cout_drain_IO_L1_out_wrapper386_U0_fifo_cout_drain_out_V_V_write_pass_0_in;
  wire [63:0] cout_drain_IO_L1_out_wrapper404_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_2_10_V_V_full_n_pass_0_in;
  wire cout_drain_IO_L1_out_wrapper404_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper283_U0_fifo_cin_out_V_V_din_pass_0_out;
  wire fifo_cin_PE_12_1_V_V_full_n_pass_0_in;
  wire PE_wrapper283_U0_fifo_cin_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper258_U0_fifo_cin_out_V_V_din_pass_0_in;
  wire fifo_cin_PE_10_0_V_V_full_n_pass_0_out;
  wire PE_wrapper258_U0_fifo_cin_out_V_V_write_pass_0_in;
  wire [63:0] cout_drain_IO_L1_out_wrapper369_U0_fifo_cout_drain_out_V_V_din_pass_1_in;
  wire fifo_cout_drain_cout_drain_IO_L1_out_0_13_V_V_full_n_pass_1_out;
  wire cout_drain_IO_L1_out_wrapper369_U0_fifo_cout_drain_out_V_V_write_pass_1_in;
  wire [255:0] PE_wrapper270_U0_fifo_w_out_V_V_din_pass_0_out;
  wire fifo_w_PE_10_1_V_V_full_n_pass_0_in;
  wire PE_wrapper270_U0_fifo_w_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper284_U0_fifo_w_out_V_V_din_pass_0_out;
  wire fifo_w_PE_11_3_V_V_full_n_pass_0_in;
  wire PE_wrapper284_U0_fifo_w_out_V_V_write_pass_0_out;
  wire [63:0] cout_drain_IO_L1_out_wrapper390_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_1_8_V_V_full_n_pass_0_in;
  wire cout_drain_IO_L1_out_wrapper390_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  wire [31:0] PE_wrapper259_U0_fifo_cout_drain_out_V_din_pass_0_in;
  wire fifo_cout_drain_PE_9_1_V_full_n_pass_0_out;
  wire PE_wrapper259_U0_fifo_cout_drain_out_V_write_pass_0_in;
  wire [255:0] PE_wrapper272_U0_fifo_w_out_V_V_din_pass_0_out;
  wire fifo_w_PE_10_3_V_V_full_n_pass_0_in;
  wire PE_wrapper272_U0_fifo_w_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper284_U0_fifo_cin_out_V_V_din_pass_0_out;
  wire fifo_cin_PE_12_2_V_V_full_n_pass_0_in;
  wire PE_wrapper284_U0_fifo_cin_out_V_V_write_pass_0_out;
  wire [31:0] PE_wrapper271_U0_fifo_cout_drain_out_V_din_pass_0_in;
  wire fifo_cout_drain_PE_10_1_V_full_n_pass_0_out;
  wire PE_wrapper271_U0_fifo_cout_drain_out_V_write_pass_0_in;
  wire ap_start_Boundary_X0Y2_To_X2Y2_in;
  wire ap_rst_n_Boundary_X0Y2_To_X2Y2_in;
  wire ap_done_Boundary_X0Y2_To_X2Y2_out;
  wire ap_start_Boundary_X0Y4_To_X2Y4_out;
  wire ap_rst_n_Boundary_X0Y4_To_X2Y4_out;
  wire ap_done_Boundary_X0Y4_To_X2Y4_in;
  wire [255:0] PE_wrapper212_U0_fifo_cin_out_V_V_din_pass_1_in;
  wire [255:0] PE_wrapper212_U0_fifo_cin_out_V_V_din_pass_2_out;
  wire fifo_cin_PE_6_2_V_V_full_n_pass_1_out;
  wire fifo_cin_PE_6_2_V_V_full_n_pass_2_in;
  wire PE_wrapper212_U0_fifo_cin_out_V_V_write_pass_1_in;
  wire PE_wrapper212_U0_fifo_cin_out_V_V_write_pass_2_out;
  wire [255:0] PE_wrapper213_U0_fifo_cin_out_V_V_din_pass_1_in;
  wire [255:0] PE_wrapper213_U0_fifo_cin_out_V_V_din_pass_2_out;
  wire fifo_cin_PE_6_3_V_V_full_n_pass_1_out;
  wire fifo_cin_PE_6_3_V_V_full_n_pass_2_in;
  wire PE_wrapper213_U0_fifo_cin_out_V_V_write_pass_1_in;
  wire PE_wrapper213_U0_fifo_cin_out_V_V_write_pass_2_out;
  wire [63:0] cout_drain_IO_L1_out_wrapper374_U0_fifo_cout_drain_out_V_V_din_pass_0_in;
  wire [63:0] cout_drain_IO_L1_out_wrapper374_U0_fifo_cout_drain_out_V_V_din_pass_1_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_0_8_V_V_full_n_pass_0_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_0_8_V_V_full_n_pass_1_in;
  wire cout_drain_IO_L1_out_wrapper374_U0_fifo_cout_drain_out_V_V_write_pass_0_in;
  wire cout_drain_IO_L1_out_wrapper374_U0_fifo_cout_drain_out_V_V_write_pass_1_out;
  wire [255:0] w_IO_L2_in140_U0_fifo_w_out_V_V_din_pass_2_in;
  wire fifo_w_w_IO_L2_in_6_V_V_full_n_pass_2_out;
  wire w_IO_L2_in140_U0_fifo_w_out_V_V_write_pass_2_in;
  wire [255:0] PE_wrapper260_U0_fifo_cin_out_V_V_din_pass_0_out;
  wire fifo_cin_PE_10_2_V_V_full_n_pass_0_in;
  wire PE_wrapper260_U0_fifo_cin_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper224_U0_fifo_cin_out_V_V_din_pass_0_in;
  wire fifo_cin_PE_7_2_V_V_full_n_pass_0_out;
  wire PE_wrapper224_U0_fifo_cin_out_V_V_write_pass_0_in;
  wire [255:0] PE_wrapper261_U0_fifo_w_out_V_V_din_pass_0_out;
  wire fifo_w_PE_9_4_V_V_full_n_pass_0_in;
  wire PE_wrapper261_U0_fifo_w_out_V_V_write_pass_0_out;
  wire [31:0] PE_wrapper235_U0_fifo_cout_drain_out_V_din_pass_0_in;
  wire fifo_cout_drain_PE_7_1_V_full_n_pass_0_out;
  wire PE_wrapper235_U0_fifo_cout_drain_out_V_write_pass_0_in;
  wire [31:0] PE_wrapper225_U0_fifo_cout_drain_out_V_din_pass_0_in;
  wire fifo_cout_drain_PE_6_3_V_full_n_pass_0_out;
  wire PE_wrapper225_U0_fifo_cout_drain_out_V_write_pass_0_in;
  wire [255:0] w_IO_L2_in141_U0_fifo_w_out_V_V_din_pass_0_out;
  wire fifo_w_w_IO_L2_in_7_V_V_full_n_pass_0_in;
  wire w_IO_L2_in141_U0_fifo_w_out_V_V_write_pass_0_out;
  wire [31:0] PE_wrapper222_U0_fifo_cout_drain_out_V_din_pass_0_in;
  wire fifo_cout_drain_PE_6_0_V_full_n_pass_0_out;
  wire PE_wrapper222_U0_fifo_cout_drain_out_V_write_pass_0_in;
  wire [255:0] PE_wrapper247_U0_fifo_w_out_V_V_din_pass_0_in;
  wire fifo_w_PE_8_2_V_V_full_n_pass_0_out;
  wire PE_wrapper247_U0_fifo_w_out_V_V_write_pass_0_in;
  wire [63:0] cout_drain_IO_L1_out_wrapper424_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_3_6_V_V_full_n_pass_0_in;
  wire cout_drain_IO_L1_out_wrapper424_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper211_U0_fifo_cin_out_V_V_din_pass_1_in;
  wire fifo_cin_PE_6_1_V_V_full_n_pass_1_out;
  wire PE_wrapper211_U0_fifo_cin_out_V_V_write_pass_1_in;
  wire [63:0] cout_drain_IO_L1_out_wrapper421_U0_fifo_cout_drain_out_V_V_din_pass_0_in;
  wire fifo_cout_drain_cout_drain_IO_L1_out_3_9_V_V_full_n_pass_0_out;
  wire cout_drain_IO_L1_out_wrapper421_U0_fifo_cout_drain_out_V_V_write_pass_0_in;
  wire [255:0] w_IO_L2_in141_U0_fifo_w_local_out_V_V_din_pass_0_out;
  wire fifo_w_PE_6_0_V_V_full_n_pass_0_in;
  wire w_IO_L2_in141_U0_fifo_w_local_out_V_V_write_pass_0_out;
  wire [31:0] PE_wrapper261_U0_fifo_cout_drain_out_V_din_pass_0_out;
  wire fifo_cout_drain_PE_9_3_V_full_n_pass_0_in;
  wire PE_wrapper261_U0_fifo_cout_drain_out_V_write_pass_0_out;
  wire [255:0] PE_wrapper222_U0_fifo_w_out_V_V_din_pass_0_in;
  wire fifo_w_PE_6_1_V_V_full_n_pass_0_out;
  wire PE_wrapper222_U0_fifo_w_out_V_V_write_pass_0_in;
  wire [63:0] cout_drain_IO_L1_out_wrapper376_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_0_6_V_V_full_n_pass_0_in;
  wire cout_drain_IO_L1_out_wrapper376_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper236_U0_fifo_w_out_V_V_din_pass_0_out;
  wire fifo_w_PE_7_3_V_V_full_n_pass_0_in;
  wire PE_wrapper236_U0_fifo_w_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper223_U0_fifo_cin_out_V_V_din_pass_0_out;
  wire fifo_cin_PE_7_1_V_V_full_n_pass_0_in;
  wire PE_wrapper223_U0_fifo_cin_out_V_V_write_pass_0_out;
  wire [63:0] cout_drain_IO_L1_out_wrapper404_U0_fifo_cout_drain_out_V_V_din_pass_1_in;
  wire fifo_cout_drain_cout_drain_IO_L1_out_2_10_V_V_full_n_pass_1_out;
  wire cout_drain_IO_L1_out_wrapper404_U0_fifo_cout_drain_out_V_V_write_pass_1_in;
  wire [255:0] PE_wrapper249_U0_fifo_w_out_V_V_din_pass_0_out;
  wire fifo_w_PE_8_4_V_V_full_n_pass_0_in;
  wire PE_wrapper249_U0_fifo_w_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper223_U0_fifo_w_out_V_V_din_pass_0_out;
  wire fifo_w_PE_6_2_V_V_full_n_pass_0_in;
  wire PE_wrapper223_U0_fifo_w_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper259_U0_fifo_w_out_V_V_din_pass_0_in;
  wire fifo_w_PE_9_2_V_V_full_n_pass_0_out;
  wire PE_wrapper259_U0_fifo_w_out_V_V_write_pass_0_in;
  wire [63:0] cout_drain_IO_L1_out_wrapper390_U0_fifo_cout_drain_out_V_V_din_pass_1_in;
  wire fifo_cout_drain_cout_drain_IO_L1_out_1_8_V_V_full_n_pass_1_out;
  wire cout_drain_IO_L1_out_wrapper390_U0_fifo_cout_drain_out_V_V_write_pass_1_in;
  wire [255:0] PE_wrapper237_U0_fifo_cin_out_V_V_din_pass_0_in;
  wire fifo_cin_PE_8_3_V_V_full_n_pass_0_out;
  wire PE_wrapper237_U0_fifo_cin_out_V_V_write_pass_0_in;
  wire [63:0] cout_drain_IO_L1_out_wrapper408_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_2_6_V_V_full_n_pass_0_in;
  wire cout_drain_IO_L1_out_wrapper408_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  wire [31:0] PE_wrapper224_U0_fifo_cout_drain_out_V_din_pass_0_in;
  wire fifo_cout_drain_PE_6_2_V_full_n_pass_0_out;
  wire PE_wrapper224_U0_fifo_cout_drain_out_V_write_pass_0_in;
  wire [255:0] PE_wrapper235_U0_fifo_w_out_V_V_din_pass_0_in;
  wire fifo_w_PE_7_2_V_V_full_n_pass_0_out;
  wire PE_wrapper235_U0_fifo_w_out_V_V_write_pass_0_in;
  wire [255:0] PE_wrapper261_U0_fifo_cin_out_V_V_din_pass_0_out;
  wire fifo_cin_PE_10_3_V_V_full_n_pass_0_in;
  wire PE_wrapper261_U0_fifo_cin_out_V_V_write_pass_0_out;
  wire [63:0] cout_drain_IO_L1_out_wrapper375_U0_fifo_cout_drain_out_V_V_din_pass_0_in;
  wire fifo_cout_drain_cout_drain_IO_L1_out_0_7_V_V_full_n_pass_0_out;
  wire cout_drain_IO_L1_out_wrapper375_U0_fifo_cout_drain_out_V_V_write_pass_0_in;
  wire [63:0] cout_drain_IO_L1_out_wrapper392_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_1_6_V_V_full_n_pass_0_in;
  wire cout_drain_IO_L1_out_wrapper392_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  wire [31:0] PE_wrapper237_U0_fifo_cout_drain_out_V_din_pass_0_in;
  wire fifo_cout_drain_PE_7_3_V_full_n_pass_0_out;
  wire PE_wrapper237_U0_fifo_cout_drain_out_V_write_pass_0_in;
  wire ap_start_Boundary_X4Y0_To_X4Y2_in;
  wire ap_rst_n_Boundary_X4Y0_To_X4Y2_in;
  wire ap_done_Boundary_X4Y0_To_X4Y2_out;
  wire ap_start_Boundary_X2Y2_To_X4Y2_out;
  wire ap_rst_n_Boundary_X2Y2_To_X4Y2_out;
  wire ap_done_Boundary_X2Y2_To_X4Y2_in;
  wire ap_start_Boundary_X2Y0_To_X2Y2_out;
  wire ap_rst_n_Boundary_X2Y0_To_X2Y2_out;
  wire ap_done_Boundary_X2Y0_To_X2Y2_in;
  wire [255:0] w_IO_L2_in140_U0_fifo_w_out_V_V_din_pass_1_in;
  wire [255:0] w_IO_L2_in140_U0_fifo_w_out_V_V_din_pass_2_out;
  wire fifo_w_w_IO_L2_in_6_V_V_full_n_pass_1_out;
  wire fifo_w_w_IO_L2_in_6_V_V_full_n_pass_2_in;
  wire w_IO_L2_in140_U0_fifo_w_out_V_V_write_pass_1_in;
  wire w_IO_L2_in140_U0_fifo_w_out_V_V_write_pass_2_out;
  wire [63:0] cout_drain_IO_L1_out_wrapper404_U0_fifo_cout_drain_out_V_V_din_pass_0_in;
  wire [63:0] cout_drain_IO_L1_out_wrapper404_U0_fifo_cout_drain_out_V_V_din_pass_1_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_2_10_V_V_full_n_pass_0_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_2_10_V_V_full_n_pass_1_in;
  wire cout_drain_IO_L1_out_wrapper404_U0_fifo_cout_drain_out_V_V_write_pass_0_in;
  wire cout_drain_IO_L1_out_wrapper404_U0_fifo_cout_drain_out_V_V_write_pass_1_out;
  wire [63:0] cout_drain_IO_L1_out_wrapper390_U0_fifo_cout_drain_out_V_V_din_pass_0_in;
  wire [63:0] cout_drain_IO_L1_out_wrapper390_U0_fifo_cout_drain_out_V_V_din_pass_1_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_1_8_V_V_full_n_pass_0_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_1_8_V_V_full_n_pass_1_in;
  wire cout_drain_IO_L1_out_wrapper390_U0_fifo_cout_drain_out_V_V_write_pass_0_in;
  wire cout_drain_IO_L1_out_wrapper390_U0_fifo_cout_drain_out_V_V_write_pass_1_out;
  wire [255:0] PE_wrapper249_U0_fifo_w_out_V_V_din_pass_0_in;
  wire [255:0] PE_wrapper249_U0_fifo_w_out_V_V_din_pass_1_out;
  wire fifo_w_PE_8_4_V_V_full_n_pass_0_out;
  wire fifo_w_PE_8_4_V_V_full_n_pass_1_in;
  wire PE_wrapper249_U0_fifo_w_out_V_V_write_pass_0_in;
  wire PE_wrapper249_U0_fifo_w_out_V_V_write_pass_1_out;
  wire [255:0] PE_wrapper272_U0_fifo_w_out_V_V_din_pass_0_in;
  wire [255:0] PE_wrapper272_U0_fifo_w_out_V_V_din_pass_1_out;
  wire fifo_w_PE_10_3_V_V_full_n_pass_0_out;
  wire fifo_w_PE_10_3_V_V_full_n_pass_1_in;
  wire PE_wrapper272_U0_fifo_w_out_V_V_write_pass_0_in;
  wire PE_wrapper272_U0_fifo_w_out_V_V_write_pass_1_out;
  wire [255:0] PE_wrapper261_U0_fifo_cin_out_V_V_din_pass_0_in;
  wire [255:0] PE_wrapper261_U0_fifo_cin_out_V_V_din_pass_1_out;
  wire fifo_cin_PE_10_3_V_V_full_n_pass_0_out;
  wire fifo_cin_PE_10_3_V_V_full_n_pass_1_in;
  wire PE_wrapper261_U0_fifo_cin_out_V_V_write_pass_0_in;
  wire PE_wrapper261_U0_fifo_cin_out_V_V_write_pass_1_out;
  wire [255:0] PE_wrapper224_U0_fifo_cin_out_V_V_din_pass_0_out;
  wire fifo_cin_PE_7_2_V_V_full_n_pass_0_in;
  wire PE_wrapper224_U0_fifo_cin_out_V_V_write_pass_0_out;
  wire [31:0] PE_wrapper235_U0_fifo_cout_drain_out_V_din_pass_0_out;
  wire fifo_cout_drain_PE_7_1_V_full_n_pass_0_in;
  wire PE_wrapper235_U0_fifo_cout_drain_out_V_write_pass_0_out;
  wire [31:0] PE_wrapper225_U0_fifo_cout_drain_out_V_din_pass_0_out;
  wire fifo_cout_drain_PE_6_3_V_full_n_pass_0_in;
  wire PE_wrapper225_U0_fifo_cout_drain_out_V_write_pass_0_out;
  wire [255:0] w_IO_L2_in141_U0_fifo_w_out_V_V_din_pass_0_in;
  wire fifo_w_w_IO_L2_in_7_V_V_full_n_pass_0_out;
  wire w_IO_L2_in141_U0_fifo_w_out_V_V_write_pass_0_in;
  wire [255:0] PE_wrapper235_U0_fifo_cin_out_V_V_din_pass_0_out;
  wire fifo_cin_PE_8_1_V_V_full_n_pass_0_in;
  wire PE_wrapper235_U0_fifo_cin_out_V_V_write_pass_0_out;
  wire [31:0] PE_wrapper222_U0_fifo_cout_drain_out_V_din_pass_0_out;
  wire fifo_cout_drain_PE_6_0_V_full_n_pass_0_in;
  wire PE_wrapper222_U0_fifo_cout_drain_out_V_write_pass_0_out;
  wire [255:0] PE_wrapper212_U0_fifo_cin_out_V_V_din_pass_2_in;
  wire fifo_cin_PE_6_2_V_V_full_n_pass_2_out;
  wire PE_wrapper212_U0_fifo_cin_out_V_V_write_pass_2_in;
  wire [255:0] PE_wrapper225_U0_fifo_w_out_V_V_din_pass_0_out;
  wire fifo_w_PE_6_4_V_V_full_n_pass_0_in;
  wire PE_wrapper225_U0_fifo_w_out_V_V_write_pass_0_out;
  wire [63:0] cout_drain_IO_L1_out_wrapper421_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_3_9_V_V_full_n_pass_0_in;
  wire cout_drain_IO_L1_out_wrapper421_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  wire [255:0] w_IO_L2_in141_U0_fifo_w_local_out_V_V_din_pass_0_in;
  wire fifo_w_PE_6_0_V_V_full_n_pass_0_out;
  wire w_IO_L2_in141_U0_fifo_w_local_out_V_V_write_pass_0_in;
  wire [63:0] cout_drain_IO_L1_out_wrapper375_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_0_7_V_V_full_n_pass_0_in;
  wire cout_drain_IO_L1_out_wrapper375_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  wire [31:0] PE_wrapper261_U0_fifo_cout_drain_out_V_din_pass_0_in;
  wire fifo_cout_drain_PE_9_3_V_full_n_pass_0_out;
  wire PE_wrapper261_U0_fifo_cout_drain_out_V_write_pass_0_in;
  wire [255:0] PE_wrapper213_U0_fifo_cin_out_V_V_din_pass_2_in;
  wire fifo_cin_PE_6_3_V_V_full_n_pass_2_out;
  wire PE_wrapper213_U0_fifo_cin_out_V_V_write_pass_2_in;
  wire [255:0] PE_wrapper222_U0_fifo_w_out_V_V_din_pass_0_out;
  wire fifo_w_PE_6_1_V_V_full_n_pass_0_in;
  wire PE_wrapper222_U0_fifo_w_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper237_U0_fifo_w_out_V_V_din_pass_0_out;
  wire fifo_w_PE_7_4_V_V_full_n_pass_0_in;
  wire PE_wrapper237_U0_fifo_w_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper236_U0_fifo_w_out_V_V_din_pass_0_in;
  wire fifo_w_PE_7_3_V_V_full_n_pass_0_out;
  wire PE_wrapper236_U0_fifo_w_out_V_V_write_pass_0_in;
  wire [255:0] PE_wrapper223_U0_fifo_cin_out_V_V_din_pass_0_in;
  wire fifo_cin_PE_7_1_V_V_full_n_pass_0_out;
  wire PE_wrapper223_U0_fifo_cin_out_V_V_write_pass_0_in;
  wire [63:0] cout_drain_IO_L1_out_wrapper374_U0_fifo_cout_drain_out_V_V_din_pass_1_in;
  wire fifo_cout_drain_cout_drain_IO_L1_out_0_8_V_V_full_n_pass_1_out;
  wire cout_drain_IO_L1_out_wrapper374_U0_fifo_cout_drain_out_V_V_write_pass_1_in;
  wire [255:0] PE_wrapper223_U0_fifo_w_out_V_V_din_pass_0_in;
  wire fifo_w_PE_6_2_V_V_full_n_pass_0_out;
  wire PE_wrapper223_U0_fifo_w_out_V_V_write_pass_0_in;
  wire [63:0] cout_drain_IO_L1_out_wrapper420_U0_fifo_cout_drain_out_V_V_din_pass_0_in;
  wire fifo_cout_drain_cout_drain_IO_L1_out_3_10_V_V_full_n_pass_0_out;
  wire cout_drain_IO_L1_out_wrapper420_U0_fifo_cout_drain_out_V_V_write_pass_0_in;
  wire [255:0] PE_wrapper234_U0_fifo_cin_out_V_V_din_pass_0_out;
  wire fifo_cin_PE_8_0_V_V_full_n_pass_0_in;
  wire PE_wrapper234_U0_fifo_cin_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper237_U0_fifo_cin_out_V_V_din_pass_0_out;
  wire fifo_cin_PE_8_3_V_V_full_n_pass_0_in;
  wire PE_wrapper237_U0_fifo_cin_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper235_U0_fifo_w_out_V_V_din_pass_0_out;
  wire fifo_w_PE_7_2_V_V_full_n_pass_0_in;
  wire PE_wrapper235_U0_fifo_w_out_V_V_write_pass_0_out;
  wire [255:0] w_IO_L2_in142_U0_fifo_w_out_V_V_din_pass_0_out;
  wire fifo_w_w_IO_L2_in_8_V_V_full_n_pass_0_in;
  wire w_IO_L2_in142_U0_fifo_w_out_V_V_write_pass_0_out;
  wire [31:0] PE_wrapper224_U0_fifo_cout_drain_out_V_din_pass_0_out;
  wire fifo_cout_drain_PE_6_2_V_full_n_pass_0_in;
  wire PE_wrapper224_U0_fifo_cout_drain_out_V_write_pass_0_out;
  wire [255:0] PE_wrapper210_U0_fifo_cin_out_V_V_din_pass_1_in;
  wire fifo_cin_PE_6_0_V_V_full_n_pass_1_out;
  wire PE_wrapper210_U0_fifo_cin_out_V_V_write_pass_1_in;
  wire [31:0] PE_wrapper237_U0_fifo_cout_drain_out_V_din_pass_0_out;
  wire fifo_cout_drain_PE_7_3_V_full_n_pass_0_in;
  wire PE_wrapper237_U0_fifo_cout_drain_out_V_write_pass_0_out;
  wire ap_start_Boundary_X2Y2_To_X4Y2_in;
  wire ap_rst_n_Boundary_X2Y2_To_X4Y2_in;
  wire ap_done_Boundary_X2Y2_To_X4Y2_out;
  wire ap_start_Boundary_X2Y4_To_X4Y4_out;
  wire ap_rst_n_Boundary_X2Y4_To_X4Y4_out;
  wire ap_done_Boundary_X2Y4_To_X4Y4_in;
  wire [63:0] cout_drain_IO_L1_out_wrapper402_U0_fifo_cout_drain_out_V_V_din_pass_1_in;
  wire [63:0] cout_drain_IO_L1_out_wrapper402_U0_fifo_cout_drain_out_V_V_din_pass_2_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_2_12_V_V_full_n_pass_1_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_2_12_V_V_full_n_pass_2_in;
  wire cout_drain_IO_L1_out_wrapper402_U0_fifo_cout_drain_out_V_V_write_pass_1_in;
  wire cout_drain_IO_L1_out_wrapper402_U0_fifo_cout_drain_out_V_V_write_pass_2_out;
  wire [31:0] PE_wrapper294_U0_fifo_cout_drain_out_V_din_pass_0_in;
  wire [31:0] PE_wrapper294_U0_fifo_cout_drain_out_V_din_pass_1_out;
  wire fifo_cout_drain_PE_12_0_V_full_n_pass_0_out;
  wire fifo_cout_drain_PE_12_0_V_full_n_pass_1_in;
  wire PE_wrapper294_U0_fifo_cout_drain_out_V_write_pass_0_in;
  wire PE_wrapper294_U0_fifo_cout_drain_out_V_write_pass_1_out;
  wire [63:0] cout_drain_IO_L1_out_wrapper369_U0_fifo_cout_drain_out_V_V_din_pass_0_in;
  wire [63:0] cout_drain_IO_L1_out_wrapper369_U0_fifo_cout_drain_out_V_V_din_pass_1_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_0_13_V_V_full_n_pass_0_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_0_13_V_V_full_n_pass_1_in;
  wire cout_drain_IO_L1_out_wrapper369_U0_fifo_cout_drain_out_V_V_write_pass_0_in;
  wire cout_drain_IO_L1_out_wrapper369_U0_fifo_cout_drain_out_V_V_write_pass_1_out;
  wire [255:0] PE_wrapper298_U0_fifo_cin_out_V_V_din_pass_0_in;
  wire [255:0] PE_wrapper298_U0_fifo_cin_out_V_V_din_pass_1_out;
  wire fifo_cin_PE_13_4_V_V_full_n_pass_0_out;
  wire fifo_cin_PE_13_4_V_V_full_n_pass_1_in;
  wire PE_wrapper298_U0_fifo_cin_out_V_V_write_pass_0_in;
  wire PE_wrapper298_U0_fifo_cin_out_V_V_write_pass_1_out;
  wire [31:0] PE_wrapper250_U0_fifo_cout_drain_out_V_din_pass_0_in;
  wire [31:0] PE_wrapper250_U0_fifo_cout_drain_out_V_din_pass_1_out;
  wire fifo_cout_drain_PE_8_4_V_full_n_pass_0_out;
  wire fifo_cout_drain_PE_8_4_V_full_n_pass_1_in;
  wire PE_wrapper250_U0_fifo_cout_drain_out_V_write_pass_0_in;
  wire PE_wrapper250_U0_fifo_cout_drain_out_V_write_pass_1_out;
  wire [255:0] PE_wrapper282_U0_fifo_cin_out_V_V_din_pass_0_in;
  wire [255:0] PE_wrapper282_U0_fifo_cin_out_V_V_din_pass_1_out;
  wire fifo_cin_PE_12_0_V_V_full_n_pass_0_out;
  wire fifo_cin_PE_12_0_V_V_full_n_pass_1_in;
  wire PE_wrapper282_U0_fifo_cin_out_V_V_write_pass_0_in;
  wire PE_wrapper282_U0_fifo_cin_out_V_V_write_pass_1_out;
  wire [255:0] PE_wrapper237_U0_fifo_w_out_V_V_din_pass_1_in;
  wire [255:0] PE_wrapper237_U0_fifo_w_out_V_V_din_pass_2_out;
  wire fifo_w_PE_7_4_V_V_full_n_pass_1_out;
  wire fifo_w_PE_7_4_V_V_full_n_pass_2_in;
  wire PE_wrapper237_U0_fifo_w_out_V_V_write_pass_1_in;
  wire PE_wrapper237_U0_fifo_w_out_V_V_write_pass_2_out;
  wire [255:0] PE_wrapper283_U0_fifo_cin_out_V_V_din_pass_0_in;
  wire [255:0] PE_wrapper283_U0_fifo_cin_out_V_V_din_pass_1_out;
  wire fifo_cin_PE_12_1_V_V_full_n_pass_0_out;
  wire fifo_cin_PE_12_1_V_V_full_n_pass_1_in;
  wire PE_wrapper283_U0_fifo_cin_out_V_V_write_pass_0_in;
  wire PE_wrapper283_U0_fifo_cin_out_V_V_write_pass_1_out;
  wire [255:0] PE_wrapper298_U0_fifo_w_out_V_V_din_pass_0_in;
  wire [255:0] PE_wrapper298_U0_fifo_w_out_V_V_din_pass_1_out;
  wire fifo_w_PE_12_5_V_V_full_n_pass_0_out;
  wire fifo_w_PE_12_5_V_V_full_n_pass_1_in;
  wire PE_wrapper298_U0_fifo_w_out_V_V_write_pass_0_in;
  wire PE_wrapper298_U0_fifo_w_out_V_V_write_pass_1_out;
  wire [255:0] PE_wrapper322_U0_fifo_w_out_V_V_din_pass_0_in;
  wire [255:0] PE_wrapper322_U0_fifo_w_out_V_V_din_pass_1_out;
  wire fifo_w_PE_14_5_V_V_full_n_pass_0_out;
  wire fifo_w_PE_14_5_V_V_full_n_pass_1_in;
  wire PE_wrapper322_U0_fifo_w_out_V_V_write_pass_0_in;
  wire PE_wrapper322_U0_fifo_w_out_V_V_write_pass_1_out;
  wire [255:0] PE_wrapper334_U0_fifo_w_out_V_V_din_pass_0_in;
  wire [255:0] PE_wrapper334_U0_fifo_w_out_V_V_din_pass_1_out;
  wire fifo_w_PE_15_5_V_V_full_n_pass_0_out;
  wire fifo_w_PE_15_5_V_V_full_n_pass_1_in;
  wire PE_wrapper334_U0_fifo_w_out_V_V_write_pass_0_in;
  wire PE_wrapper334_U0_fifo_w_out_V_V_write_pass_1_out;
  wire [63:0] cout_drain_IO_L1_out_wrapper385_U0_fifo_cout_drain_out_V_V_din_pass_0_in;
  wire fifo_cout_drain_cout_drain_IO_L1_out_1_13_V_V_full_n_pass_0_out;
  wire cout_drain_IO_L1_out_wrapper385_U0_fifo_cout_drain_out_V_V_write_pass_0_in;
  wire [255:0] PE_wrapper309_U0_fifo_cin_out_V_V_din_pass_0_out;
  wire fifo_cin_PE_14_3_V_V_full_n_pass_0_in;
  wire PE_wrapper309_U0_fifo_cin_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper261_U0_fifo_w_out_V_V_din_pass_2_in;
  wire fifo_w_PE_9_4_V_V_full_n_pass_2_out;
  wire PE_wrapper261_U0_fifo_w_out_V_V_write_pass_2_in;
  wire [255:0] PE_wrapper333_U0_fifo_w_out_V_V_din_pass_0_out;
  wire fifo_w_PE_15_4_V_V_full_n_pass_0_in;
  wire PE_wrapper333_U0_fifo_w_out_V_V_write_pass_0_out;
  wire [63:0] cout_drain_IO_L1_out_wrapper440_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_4_6_V_V_full_n_pass_0_in;
  wire cout_drain_IO_L1_out_wrapper440_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper250_U0_fifo_cin_out_V_V_din_pass_0_in;
  wire fifo_cin_PE_9_4_V_V_full_n_pass_0_out;
  wire PE_wrapper250_U0_fifo_cin_out_V_V_write_pass_0_in;
  wire [31:0] PE_wrapper286_U0_fifo_cout_drain_out_V_din_pass_1_in;
  wire fifo_cout_drain_PE_11_4_V_full_n_pass_1_out;
  wire PE_wrapper286_U0_fifo_cout_drain_out_V_write_pass_1_in;
  wire [63:0] cout_drain_IO_L1_out_wrapper439_U0_fifo_cout_drain_out_V_V_din_pass_0_in;
  wire fifo_cout_drain_cout_drain_IO_L1_out_4_7_V_V_full_n_pass_0_out;
  wire cout_drain_IO_L1_out_wrapper439_U0_fifo_cout_drain_out_V_V_write_pass_0_in;
  wire [31:0] PE_wrapper306_U0_fifo_cout_drain_out_V_din_pass_0_out;
  wire fifo_cout_drain_PE_13_0_V_full_n_pass_0_in;
  wire PE_wrapper306_U0_fifo_cout_drain_out_V_write_pass_0_out;
  wire [255:0] PE_wrapper295_U0_fifo_w_out_V_V_din_pass_0_in;
  wire fifo_w_PE_12_2_V_V_full_n_pass_0_out;
  wire PE_wrapper295_U0_fifo_w_out_V_V_write_pass_0_in;
  wire [31:0] PE_wrapper226_U0_fifo_cout_drain_out_V_din_pass_1_in;
  wire fifo_cout_drain_PE_6_4_V_full_n_pass_1_out;
  wire PE_wrapper226_U0_fifo_cout_drain_out_V_write_pass_1_in;
  wire [255:0] PE_wrapper320_U0_fifo_cin_out_V_V_din_pass_1_in;
  wire fifo_cin_PE_15_2_V_V_full_n_pass_1_out;
  wire PE_wrapper320_U0_fifo_cin_out_V_V_write_pass_1_in;
  wire [255:0] PE_wrapper309_U0_fifo_w_out_V_V_din_pass_0_out;
  wire fifo_w_PE_13_4_V_V_full_n_pass_0_in;
  wire PE_wrapper309_U0_fifo_w_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper331_U0_fifo_w_out_V_V_din_pass_0_in;
  wire fifo_w_PE_15_2_V_V_full_n_pass_0_out;
  wire PE_wrapper331_U0_fifo_w_out_V_V_write_pass_0_in;
  wire [63:0] cout_drain_IO_L1_out_wrapper418_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_3_12_V_V_full_n_pass_0_in;
  wire cout_drain_IO_L1_out_wrapper418_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  wire [63:0] cout_drain_IO_L1_out_wrapper417_U0_fifo_cout_drain_out_V_V_din_pass_0_in;
  wire fifo_cout_drain_cout_drain_IO_L1_out_3_13_V_V_full_n_pass_0_out;
  wire cout_drain_IO_L1_out_wrapper417_U0_fifo_cout_drain_out_V_V_write_pass_0_in;
  wire [255:0] w_IO_L2_in147_U0_fifo_w_out_V_V_din_pass_0_out;
  wire fifo_w_w_IO_L2_in_13_V_V_full_n_pass_0_in;
  wire w_IO_L2_in147_U0_fifo_w_out_V_V_write_pass_0_out;
  wire [255:0] w_IO_L2_in146_U0_fifo_w_out_V_V_din_pass_0_in;
  wire fifo_w_w_IO_L2_in_12_V_V_full_n_pass_0_out;
  wire w_IO_L2_in146_U0_fifo_w_out_V_V_write_pass_0_in;
  wire [255:0] PE_wrapper297_U0_fifo_cin_out_V_V_din_pass_0_in;
  wire fifo_cin_PE_13_3_V_V_full_n_pass_0_out;
  wire PE_wrapper297_U0_fifo_cin_out_V_V_write_pass_0_in;
  wire [255:0] PE_wrapper285_U0_fifo_w_out_V_V_din_pass_0_out;
  wire fifo_w_PE_11_4_V_V_full_n_pass_0_in;
  wire PE_wrapper285_U0_fifo_w_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper306_U0_fifo_w_out_V_V_din_pass_0_out;
  wire fifo_w_PE_13_1_V_V_full_n_pass_0_in;
  wire PE_wrapper306_U0_fifo_w_out_V_V_write_pass_0_out;
  wire [31:0] PE_wrapper333_U0_fifo_cout_drain_out_V_din_pass_0_out;
  wire fifo_cout_drain_PE_15_3_V_full_n_pass_0_in;
  wire PE_wrapper333_U0_fifo_cout_drain_out_V_write_pass_0_out;
  wire [63:0] cout_drain_IO_L1_out_wrapper386_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_1_12_V_V_full_n_pass_0_in;
  wire cout_drain_IO_L1_out_wrapper386_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper262_U0_fifo_w_out_V_V_din_pass_0_out;
  wire fifo_w_PE_9_5_V_V_full_n_pass_0_in;
  wire PE_wrapper262_U0_fifo_w_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper306_U0_fifo_cin_out_V_V_din_pass_0_out;
  wire fifo_cin_PE_14_0_V_V_full_n_pass_0_in;
  wire PE_wrapper306_U0_fifo_cin_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper273_U0_fifo_cin_out_V_V_din_pass_0_in;
  wire fifo_cin_PE_11_3_V_V_full_n_pass_0_out;
  wire PE_wrapper273_U0_fifo_cin_out_V_V_write_pass_0_in;
  wire [255:0] PE_wrapper321_U0_fifo_cin_out_V_V_din_pass_1_in;
  wire fifo_cin_PE_15_3_V_V_full_n_pass_1_out;
  wire PE_wrapper321_U0_fifo_cin_out_V_V_write_pass_1_in;
  wire [31:0] PE_wrapper295_U0_fifo_cout_drain_out_V_din_pass_0_in;
  wire fifo_cout_drain_PE_12_1_V_full_n_pass_0_out;
  wire PE_wrapper295_U0_fifo_cout_drain_out_V_write_pass_0_in;
  wire [31:0] PE_wrapper285_U0_fifo_cout_drain_out_V_din_pass_0_out;
  wire fifo_cout_drain_PE_11_3_V_full_n_pass_0_in;
  wire PE_wrapper285_U0_fifo_cout_drain_out_V_write_pass_0_out;
  wire [255:0] PE_wrapper294_U0_fifo_cin_out_V_V_din_pass_0_in;
  wire fifo_cin_PE_13_0_V_V_full_n_pass_0_out;
  wire PE_wrapper294_U0_fifo_cin_out_V_V_write_pass_0_in;
  wire [255:0] w_IO_L2_in147_U0_fifo_w_local_out_V_V_din_pass_0_out;
  wire fifo_w_PE_12_0_V_V_full_n_pass_0_in;
  wire w_IO_L2_in147_U0_fifo_w_local_out_V_V_write_pass_0_out;
  wire [63:0] cout_drain_IO_L1_out_wrapper437_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_4_9_V_V_full_n_pass_0_in;
  wire cout_drain_IO_L1_out_wrapper437_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  wire [31:0] PE_wrapper297_U0_fifo_cout_drain_out_V_din_pass_0_in;
  wire fifo_cout_drain_PE_12_3_V_full_n_pass_0_out;
  wire PE_wrapper297_U0_fifo_cout_drain_out_V_write_pass_0_in;
  wire [255:0] PE_wrapper308_U0_fifo_w_out_V_V_din_pass_0_in;
  wire fifo_w_PE_13_3_V_V_full_n_pass_0_out;
  wire PE_wrapper308_U0_fifo_w_out_V_V_write_pass_0_in;
  wire [255:0] PE_wrapper296_U0_fifo_cin_out_V_V_din_pass_0_out;
  wire fifo_cin_PE_13_2_V_V_full_n_pass_0_in;
  wire PE_wrapper296_U0_fifo_cin_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper284_U0_fifo_w_out_V_V_din_pass_0_in;
  wire fifo_w_PE_11_3_V_V_full_n_pass_0_out;
  wire PE_wrapper284_U0_fifo_w_out_V_V_write_pass_0_in;
  wire [255:0] PE_wrapper296_U0_fifo_w_out_V_V_din_pass_0_out;
  wire fifo_w_PE_12_3_V_V_full_n_pass_0_in;
  wire PE_wrapper296_U0_fifo_w_out_V_V_write_pass_0_out;
  wire [31:0] PE_wrapper296_U0_fifo_cout_drain_out_V_din_pass_0_out;
  wire fifo_cout_drain_PE_12_2_V_full_n_pass_0_in;
  wire PE_wrapper296_U0_fifo_cout_drain_out_V_write_pass_0_out;
  wire [255:0] PE_wrapper262_U0_fifo_cin_out_V_V_din_pass_0_out;
  wire fifo_cin_PE_10_4_V_V_full_n_pass_0_in;
  wire PE_wrapper262_U0_fifo_cin_out_V_V_write_pass_0_out;
  wire [31:0] PE_wrapper274_U0_fifo_cout_drain_out_V_din_pass_1_in;
  wire fifo_cout_drain_PE_10_4_V_full_n_pass_1_out;
  wire PE_wrapper274_U0_fifo_cout_drain_out_V_write_pass_1_in;
  wire [255:0] w_IO_L2_in148_U0_fifo_w_local_out_V_V_din_pass_0_in;
  wire fifo_w_PE_13_0_V_V_full_n_pass_0_out;
  wire w_IO_L2_in148_U0_fifo_w_local_out_V_V_write_pass_0_in;
  wire [63:0] cout_drain_IO_L1_out_boundary_wrapper399_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_2_15_V_V_full_n_pass_0_in;
  wire cout_drain_IO_L1_out_boundary_wrapper399_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper284_U0_fifo_cin_out_V_V_din_pass_0_in;
  wire fifo_cin_PE_12_2_V_V_full_n_pass_0_out;
  wire PE_wrapper284_U0_fifo_cin_out_V_V_write_pass_0_in;
  wire [63:0] cout_drain_IO_L1_out_wrapper434_U0_fifo_cout_drain_out_V_V_din_pass_1_in;
  wire fifo_cout_drain_cout_drain_IO_L1_out_4_12_V_V_full_n_pass_1_out;
  wire cout_drain_IO_L1_out_wrapper434_U0_fifo_cout_drain_out_V_V_write_pass_1_in;
  wire [255:0] PE_wrapper285_U0_fifo_cin_out_V_V_din_pass_0_out;
  wire fifo_cin_PE_12_3_V_V_full_n_pass_0_in;
  wire PE_wrapper285_U0_fifo_cin_out_V_V_write_pass_0_out;
  wire [31:0] PE_wrapper309_U0_fifo_cout_drain_out_V_din_pass_0_out;
  wire fifo_cout_drain_PE_13_3_V_full_n_pass_0_in;
  wire PE_wrapper309_U0_fifo_cout_drain_out_V_write_pass_0_out;
  wire ap_start_Boundary_X0Y4_To_X2Y4_in;
  wire ap_rst_n_Boundary_X0Y4_To_X2Y4_in;
  wire ap_done_Boundary_X0Y4_To_X2Y4_out;
  wire ap_start_Boundary_X0Y6_To_X2Y6_out;
  wire ap_rst_n_Boundary_X0Y6_To_X2Y6_out;
  wire ap_done_Boundary_X0Y6_To_X2Y6_in;
  wire [63:0] cout_drain_IO_L1_out_wrapper402_U0_fifo_cout_drain_out_V_V_din_pass_0_in;
  wire [63:0] cout_drain_IO_L1_out_wrapper402_U0_fifo_cout_drain_out_V_V_din_pass_1_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_2_12_V_V_full_n_pass_0_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_2_12_V_V_full_n_pass_1_in;
  wire cout_drain_IO_L1_out_wrapper402_U0_fifo_cout_drain_out_V_V_write_pass_0_in;
  wire cout_drain_IO_L1_out_wrapper402_U0_fifo_cout_drain_out_V_V_write_pass_1_out;
  wire [31:0] PE_wrapper286_U0_fifo_cout_drain_out_V_din_pass_0_in;
  wire [31:0] PE_wrapper286_U0_fifo_cout_drain_out_V_din_pass_1_out;
  wire fifo_cout_drain_PE_11_4_V_full_n_pass_0_out;
  wire fifo_cout_drain_PE_11_4_V_full_n_pass_1_in;
  wire PE_wrapper286_U0_fifo_cout_drain_out_V_write_pass_0_in;
  wire PE_wrapper286_U0_fifo_cout_drain_out_V_write_pass_1_out;
  wire [31:0] PE_wrapper226_U0_fifo_cout_drain_out_V_din_pass_0_in;
  wire [31:0] PE_wrapper226_U0_fifo_cout_drain_out_V_din_pass_1_out;
  wire fifo_cout_drain_PE_6_4_V_full_n_pass_0_out;
  wire fifo_cout_drain_PE_6_4_V_full_n_pass_1_in;
  wire PE_wrapper226_U0_fifo_cout_drain_out_V_write_pass_0_in;
  wire PE_wrapper226_U0_fifo_cout_drain_out_V_write_pass_1_out;
  wire [255:0] PE_wrapper320_U0_fifo_cin_out_V_V_din_pass_0_in;
  wire [255:0] PE_wrapper320_U0_fifo_cin_out_V_V_din_pass_1_out;
  wire fifo_cin_PE_15_2_V_V_full_n_pass_0_out;
  wire fifo_cin_PE_15_2_V_V_full_n_pass_1_in;
  wire PE_wrapper320_U0_fifo_cin_out_V_V_write_pass_0_in;
  wire PE_wrapper320_U0_fifo_cin_out_V_V_write_pass_1_out;
  wire [255:0] PE_wrapper321_U0_fifo_cin_out_V_V_din_pass_0_in;
  wire [255:0] PE_wrapper321_U0_fifo_cin_out_V_V_din_pass_1_out;
  wire fifo_cin_PE_15_3_V_V_full_n_pass_0_out;
  wire fifo_cin_PE_15_3_V_V_full_n_pass_1_in;
  wire PE_wrapper321_U0_fifo_cin_out_V_V_write_pass_0_in;
  wire PE_wrapper321_U0_fifo_cin_out_V_V_write_pass_1_out;
  wire [31:0] PE_wrapper274_U0_fifo_cout_drain_out_V_din_pass_0_in;
  wire [31:0] PE_wrapper274_U0_fifo_cout_drain_out_V_din_pass_1_out;
  wire fifo_cout_drain_PE_10_4_V_full_n_pass_0_out;
  wire fifo_cout_drain_PE_10_4_V_full_n_pass_1_in;
  wire PE_wrapper274_U0_fifo_cout_drain_out_V_write_pass_0_in;
  wire PE_wrapper274_U0_fifo_cout_drain_out_V_write_pass_1_out;
  wire [63:0] cout_drain_IO_L1_out_wrapper434_U0_fifo_cout_drain_out_V_V_din_pass_0_in;
  wire [63:0] cout_drain_IO_L1_out_wrapper434_U0_fifo_cout_drain_out_V_V_din_pass_1_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_4_12_V_V_full_n_pass_0_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_4_12_V_V_full_n_pass_1_in;
  wire cout_drain_IO_L1_out_wrapper434_U0_fifo_cout_drain_out_V_V_write_pass_0_in;
  wire cout_drain_IO_L1_out_wrapper434_U0_fifo_cout_drain_out_V_V_write_pass_1_out;
  wire [255:0] PE_wrapper262_U0_fifo_w_out_V_V_din_pass_0_in;
  wire [255:0] PE_wrapper262_U0_fifo_w_out_V_V_din_pass_1_out;
  wire fifo_w_PE_9_5_V_V_full_n_pass_0_out;
  wire fifo_w_PE_9_5_V_V_full_n_pass_1_in;
  wire PE_wrapper262_U0_fifo_w_out_V_V_write_pass_0_in;
  wire PE_wrapper262_U0_fifo_w_out_V_V_write_pass_1_out;
  wire [255:0] PE_wrapper298_U0_fifo_w_out_V_V_din_pass_1_in;
  wire [255:0] PE_wrapper298_U0_fifo_w_out_V_V_din_pass_2_out;
  wire fifo_w_PE_12_5_V_V_full_n_pass_1_out;
  wire fifo_w_PE_12_5_V_V_full_n_pass_2_in;
  wire PE_wrapper298_U0_fifo_w_out_V_V_write_pass_1_in;
  wire PE_wrapper298_U0_fifo_w_out_V_V_write_pass_2_out;
  wire [255:0] PE_wrapper322_U0_fifo_w_out_V_V_din_pass_1_in;
  wire [255:0] PE_wrapper322_U0_fifo_w_out_V_V_din_pass_2_out;
  wire fifo_w_PE_14_5_V_V_full_n_pass_1_out;
  wire fifo_w_PE_14_5_V_V_full_n_pass_2_in;
  wire PE_wrapper322_U0_fifo_w_out_V_V_write_pass_1_in;
  wire PE_wrapper322_U0_fifo_w_out_V_V_write_pass_2_out;
  wire [255:0] PE_wrapper334_U0_fifo_w_out_V_V_din_pass_1_in;
  wire [255:0] PE_wrapper334_U0_fifo_w_out_V_V_din_pass_2_out;
  wire fifo_w_PE_15_5_V_V_full_n_pass_1_out;
  wire fifo_w_PE_15_5_V_V_full_n_pass_2_in;
  wire PE_wrapper334_U0_fifo_w_out_V_V_write_pass_1_in;
  wire PE_wrapper334_U0_fifo_w_out_V_V_write_pass_2_out;
  wire [63:0] cout_drain_IO_L1_out_wrapper385_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_1_13_V_V_full_n_pass_0_in;
  wire cout_drain_IO_L1_out_wrapper385_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper298_U0_fifo_cin_out_V_V_din_pass_1_in;
  wire fifo_cin_PE_13_4_V_V_full_n_pass_1_out;
  wire PE_wrapper298_U0_fifo_cin_out_V_V_write_pass_1_in;
  wire [31:0] PE_wrapper250_U0_fifo_cout_drain_out_V_din_pass_1_in;
  wire fifo_cout_drain_PE_8_4_V_full_n_pass_1_out;
  wire PE_wrapper250_U0_fifo_cout_drain_out_V_write_pass_1_in;
  wire [255:0] PE_wrapper310_U0_fifo_w_out_V_V_din_pass_0_out;
  wire fifo_w_PE_13_5_V_V_full_n_pass_0_in;
  wire PE_wrapper310_U0_fifo_w_out_V_V_write_pass_0_out;
  wire [63:0] cout_drain_IO_L1_out_wrapper439_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_4_7_V_V_full_n_pass_0_in;
  wire cout_drain_IO_L1_out_wrapper439_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  wire [31:0] PE_wrapper310_U0_fifo_cout_drain_out_V_din_pass_0_out;
  wire fifo_cout_drain_PE_13_4_V_full_n_pass_0_in;
  wire PE_wrapper310_U0_fifo_cout_drain_out_V_write_pass_0_out;
  wire [255:0] PE_wrapper295_U0_fifo_w_out_V_V_din_pass_0_out;
  wire fifo_w_PE_12_2_V_V_full_n_pass_0_in;
  wire PE_wrapper295_U0_fifo_w_out_V_V_write_pass_0_out;
  wire [255:0] w_IO_L2_in148_U0_fifo_w_out_V_V_din_pass_0_out;
  wire fifo_w_w_IO_L2_in_14_V_V_full_n_pass_0_in;
  wire w_IO_L2_in148_U0_fifo_w_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper309_U0_fifo_w_out_V_V_din_pass_0_in;
  wire fifo_w_PE_13_4_V_V_full_n_pass_0_out;
  wire PE_wrapper309_U0_fifo_w_out_V_V_write_pass_0_in;
  wire [63:0] cout_drain_IO_L1_out_wrapper417_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_3_13_V_V_full_n_pass_0_in;
  wire cout_drain_IO_L1_out_wrapper417_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  wire [31:0] PE_wrapper308_U0_fifo_cout_drain_out_V_din_pass_0_out;
  wire fifo_cout_drain_PE_13_2_V_full_n_pass_0_in;
  wire PE_wrapper308_U0_fifo_cout_drain_out_V_write_pass_0_out;
  wire [255:0] w_IO_L2_in147_U0_fifo_w_out_V_V_din_pass_0_in;
  wire fifo_w_w_IO_L2_in_13_V_V_full_n_pass_0_out;
  wire w_IO_L2_in147_U0_fifo_w_out_V_V_write_pass_0_in;
  wire [255:0] PE_wrapper282_U0_fifo_cin_out_V_V_din_pass_1_in;
  wire fifo_cin_PE_12_0_V_V_full_n_pass_1_out;
  wire PE_wrapper282_U0_fifo_cin_out_V_V_write_pass_1_in;
  wire [63:0] cout_drain_IO_L1_out_wrapper416_U0_fifo_cout_drain_out_V_V_din_pass_0_in;
  wire fifo_cout_drain_cout_drain_IO_L1_out_3_14_V_V_full_n_pass_0_out;
  wire cout_drain_IO_L1_out_wrapper416_U0_fifo_cout_drain_out_V_V_write_pass_0_in;
  wire [255:0] PE_wrapper297_U0_fifo_cin_out_V_V_din_pass_0_out;
  wire fifo_cin_PE_13_3_V_V_full_n_pass_0_in;
  wire PE_wrapper297_U0_fifo_cin_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper306_U0_fifo_w_out_V_V_din_pass_0_in;
  wire fifo_w_PE_13_1_V_V_full_n_pass_0_out;
  wire PE_wrapper306_U0_fifo_w_out_V_V_write_pass_0_in;
  wire [255:0] PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0_out;
  wire fifo_cin_PE_8_4_V_V_full_n_pass_0_in;
  wire PE_wrapper238_U0_fifo_cin_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0_out;
  wire fifo_w_PE_12_4_V_V_full_n_pass_0_in;
  wire PE_wrapper297_U0_fifo_w_out_V_V_write_pass_0_out;
  wire [31:0] PE_wrapper294_U0_fifo_cout_drain_out_V_din_pass_0_out;
  wire fifo_cout_drain_PE_12_0_V_full_n_pass_0_in;
  wire PE_wrapper294_U0_fifo_cout_drain_out_V_write_pass_0_out;
  wire [255:0] PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0_out;
  wire fifo_cin_PE_14_4_V_V_full_n_pass_0_in;
  wire PE_wrapper310_U0_fifo_cin_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0_out;
  wire fifo_cin_PE_14_1_V_V_full_n_pass_0_in;
  wire PE_wrapper307_U0_fifo_cin_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper237_U0_fifo_w_out_V_V_din_pass_2_in;
  wire fifo_w_PE_7_4_V_V_full_n_pass_2_out;
  wire PE_wrapper237_U0_fifo_w_out_V_V_write_pass_2_in;
  wire [255:0] PE_wrapper283_U0_fifo_cin_out_V_V_din_pass_1_in;
  wire fifo_cin_PE_12_1_V_V_full_n_pass_1_out;
  wire PE_wrapper283_U0_fifo_cin_out_V_V_write_pass_1_in;
  wire [31:0] PE_wrapper295_U0_fifo_cout_drain_out_V_din_pass_0_out;
  wire fifo_cout_drain_PE_12_1_V_full_n_pass_0_in;
  wire PE_wrapper295_U0_fifo_cout_drain_out_V_write_pass_0_out;
  wire [255:0] PE_wrapper294_U0_fifo_cin_out_V_V_din_pass_0_out;
  wire fifo_cin_PE_13_0_V_V_full_n_pass_0_in;
  wire PE_wrapper294_U0_fifo_cin_out_V_V_write_pass_0_out;
  wire [255:0] w_IO_L2_in147_U0_fifo_w_local_out_V_V_din_pass_0_in;
  wire fifo_w_PE_12_0_V_V_full_n_pass_0_out;
  wire w_IO_L2_in147_U0_fifo_w_local_out_V_V_write_pass_0_in;
  wire [63:0] cout_drain_IO_L1_out_wrapper437_U0_fifo_cout_drain_out_V_V_din_pass_0_in;
  wire fifo_cout_drain_cout_drain_IO_L1_out_4_9_V_V_full_n_pass_0_out;
  wire cout_drain_IO_L1_out_wrapper437_U0_fifo_cout_drain_out_V_V_write_pass_0_in;
  wire [31:0] PE_wrapper297_U0_fifo_cout_drain_out_V_din_pass_0_out;
  wire fifo_cout_drain_PE_12_3_V_full_n_pass_0_in;
  wire PE_wrapper297_U0_fifo_cout_drain_out_V_write_pass_0_out;
  wire [255:0] PE_wrapper308_U0_fifo_cin_out_V_V_din_pass_0_out;
  wire fifo_cin_PE_14_2_V_V_full_n_pass_0_in;
  wire PE_wrapper308_U0_fifo_cin_out_V_V_write_pass_0_out;
  wire [63:0] cout_drain_IO_L1_out_wrapper384_U0_fifo_cout_drain_out_V_V_din_pass_0_in;
  wire fifo_cout_drain_cout_drain_IO_L1_out_1_14_V_V_full_n_pass_0_out;
  wire cout_drain_IO_L1_out_wrapper384_U0_fifo_cout_drain_out_V_V_write_pass_0_in;
  wire [255:0] PE_wrapper308_U0_fifo_w_out_V_V_din_pass_0_out;
  wire fifo_w_PE_13_3_V_V_full_n_pass_0_in;
  wire PE_wrapper308_U0_fifo_w_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper296_U0_fifo_cin_out_V_V_din_pass_0_in;
  wire fifo_cin_PE_13_2_V_V_full_n_pass_0_out;
  wire PE_wrapper296_U0_fifo_cin_out_V_V_write_pass_0_in;
  wire [255:0] PE_wrapper296_U0_fifo_w_out_V_V_din_pass_0_in;
  wire fifo_w_PE_12_3_V_V_full_n_pass_0_out;
  wire PE_wrapper296_U0_fifo_w_out_V_V_write_pass_0_in;
  wire [255:0] PE_wrapper226_U0_fifo_cin_out_V_V_din_pass_0_in;
  wire fifo_cin_PE_7_4_V_V_full_n_pass_0_out;
  wire PE_wrapper226_U0_fifo_cin_out_V_V_write_pass_0_in;
  wire [255:0] w_IO_L2_in148_U0_fifo_w_local_out_V_V_din_pass_0_out;
  wire fifo_w_PE_13_0_V_V_full_n_pass_0_in;
  wire w_IO_L2_in148_U0_fifo_w_local_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0_out;
  wire fifo_w_PE_7_5_V_V_full_n_pass_0_in;
  wire PE_wrapper238_U0_fifo_w_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper285_U0_fifo_cin_out_V_V_din_pass_0_in;
  wire fifo_cin_PE_12_3_V_V_full_n_pass_0_out;
  wire PE_wrapper285_U0_fifo_cin_out_V_V_write_pass_0_in;
  wire [31:0] PE_wrapper309_U0_fifo_cout_drain_out_V_din_pass_0_in;
  wire fifo_cout_drain_PE_13_3_V_full_n_pass_0_out;
  wire PE_wrapper309_U0_fifo_cout_drain_out_V_write_pass_0_in;
  wire ap_start_Boundary_X0Y6_To_X2Y6_in;
  wire ap_rst_n_Boundary_X0Y6_To_X2Y6_in;
  wire ap_done_Boundary_X0Y6_To_X2Y6_out;
  wire ap_start_Boundary_X0Y8_To_X2Y8_out;
  wire ap_rst_n_Boundary_X0Y8_To_X2Y8_out;
  wire ap_done_Boundary_X0Y8_To_X2Y8_in;
  wire [255:0] PE_wrapper309_U0_fifo_cin_out_V_V_din_pass_0_in;
  wire [255:0] PE_wrapper309_U0_fifo_cin_out_V_V_din_pass_1_out;
  wire fifo_cin_PE_14_3_V_V_full_n_pass_0_out;
  wire fifo_cin_PE_14_3_V_V_full_n_pass_1_in;
  wire PE_wrapper309_U0_fifo_cin_out_V_V_write_pass_0_in;
  wire PE_wrapper309_U0_fifo_cin_out_V_V_write_pass_1_out;
  wire [255:0] PE_wrapper214_U0_fifo_cin_out_V_V_din_pass_0_in;
  wire [255:0] PE_wrapper214_U0_fifo_cin_out_V_V_din_pass_1_out;
  wire fifo_cin_PE_6_4_V_V_full_n_pass_0_out;
  wire fifo_cin_PE_6_4_V_V_full_n_pass_1_in;
  wire PE_wrapper214_U0_fifo_cin_out_V_V_write_pass_0_in;
  wire PE_wrapper214_U0_fifo_cin_out_V_V_write_pass_1_out;
  wire [63:0] cout_drain_IO_L1_out_wrapper418_U0_fifo_cout_drain_out_V_V_din_pass_0_in;
  wire [63:0] cout_drain_IO_L1_out_wrapper418_U0_fifo_cout_drain_out_V_V_din_pass_1_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_3_12_V_V_full_n_pass_0_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_3_12_V_V_full_n_pass_1_in;
  wire cout_drain_IO_L1_out_wrapper418_U0_fifo_cout_drain_out_V_V_write_pass_0_in;
  wire cout_drain_IO_L1_out_wrapper418_U0_fifo_cout_drain_out_V_V_write_pass_1_out;
  wire [255:0] PE_wrapper225_U0_fifo_w_out_V_V_din_pass_0_in;
  wire [255:0] PE_wrapper225_U0_fifo_w_out_V_V_din_pass_1_out;
  wire fifo_w_PE_6_4_V_V_full_n_pass_0_out;
  wire fifo_w_PE_6_4_V_V_full_n_pass_1_in;
  wire PE_wrapper225_U0_fifo_w_out_V_V_write_pass_0_in;
  wire PE_wrapper225_U0_fifo_w_out_V_V_write_pass_1_out;
  wire [255:0] PE_wrapper285_U0_fifo_w_out_V_V_din_pass_0_in;
  wire [255:0] PE_wrapper285_U0_fifo_w_out_V_V_din_pass_1_out;
  wire fifo_w_PE_11_4_V_V_full_n_pass_0_out;
  wire fifo_w_PE_11_4_V_V_full_n_pass_1_in;
  wire PE_wrapper285_U0_fifo_w_out_V_V_write_pass_0_in;
  wire PE_wrapper285_U0_fifo_w_out_V_V_write_pass_1_out;
  wire [255:0] PE_wrapper306_U0_fifo_cin_out_V_V_din_pass_0_in;
  wire [255:0] PE_wrapper306_U0_fifo_cin_out_V_V_din_pass_1_out;
  wire fifo_cin_PE_14_0_V_V_full_n_pass_0_out;
  wire fifo_cin_PE_14_0_V_V_full_n_pass_1_in;
  wire PE_wrapper306_U0_fifo_cin_out_V_V_write_pass_0_in;
  wire PE_wrapper306_U0_fifo_cin_out_V_V_write_pass_1_out;
  wire [31:0] PE_wrapper285_U0_fifo_cout_drain_out_V_din_pass_0_in;
  wire [31:0] PE_wrapper285_U0_fifo_cout_drain_out_V_din_pass_1_out;
  wire fifo_cout_drain_PE_11_3_V_full_n_pass_0_out;
  wire fifo_cout_drain_PE_11_3_V_full_n_pass_1_in;
  wire PE_wrapper285_U0_fifo_cout_drain_out_V_write_pass_0_in;
  wire PE_wrapper285_U0_fifo_cout_drain_out_V_write_pass_1_out;
  wire [255:0] PE_wrapper262_U0_fifo_cin_out_V_V_din_pass_0_in;
  wire [255:0] PE_wrapper262_U0_fifo_cin_out_V_V_din_pass_1_out;
  wire fifo_cin_PE_10_4_V_V_full_n_pass_0_out;
  wire fifo_cin_PE_10_4_V_V_full_n_pass_1_in;
  wire PE_wrapper262_U0_fifo_cin_out_V_V_write_pass_0_in;
  wire PE_wrapper262_U0_fifo_cin_out_V_V_write_pass_1_out;
  wire [31:0] PE_wrapper296_U0_fifo_cout_drain_out_V_din_pass_0_in;
  wire [31:0] PE_wrapper296_U0_fifo_cout_drain_out_V_din_pass_1_out;
  wire fifo_cout_drain_PE_12_2_V_full_n_pass_0_out;
  wire fifo_cout_drain_PE_12_2_V_full_n_pass_1_in;
  wire PE_wrapper296_U0_fifo_cout_drain_out_V_write_pass_0_in;
  wire PE_wrapper296_U0_fifo_cout_drain_out_V_write_pass_1_out;
  wire [63:0] cout_drain_IO_L1_out_wrapper440_U0_fifo_cout_drain_out_V_V_din_pass_0_in;
  wire [63:0] cout_drain_IO_L1_out_wrapper440_U0_fifo_cout_drain_out_V_V_din_pass_1_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_4_6_V_V_full_n_pass_0_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_4_6_V_V_full_n_pass_1_in;
  wire cout_drain_IO_L1_out_wrapper440_U0_fifo_cout_drain_out_V_V_write_pass_0_in;
  wire cout_drain_IO_L1_out_wrapper440_U0_fifo_cout_drain_out_V_V_write_pass_1_out;
  wire [31:0] PE_wrapper320_U0_fifo_cout_drain_out_V_din_pass_0_in;
  wire fifo_cout_drain_PE_14_2_V_full_n_pass_0_out;
  wire PE_wrapper320_U0_fifo_cout_drain_out_V_write_pass_0_in;
  wire [63:0] cout_drain_IO_L1_out_wrapper433_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_4_13_V_V_full_n_pass_0_in;
  wire cout_drain_IO_L1_out_wrapper433_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper333_U0_fifo_w_out_V_V_din_pass_0_in;
  wire fifo_w_PE_15_4_V_V_full_n_pass_0_out;
  wire PE_wrapper333_U0_fifo_w_out_V_V_write_pass_0_in;
  wire [255:0] w_IO_L2_in149_U0_fifo_w_out_V_V_din_pass_0_in;
  wire fifo_w_w_IO_L2_in_15_V_V_full_n_pass_0_out;
  wire w_IO_L2_in149_U0_fifo_w_out_V_V_write_pass_0_in;
  wire [255:0] PE_wrapper250_U0_fifo_cin_out_V_V_din_pass_0_out;
  wire fifo_cin_PE_9_4_V_V_full_n_pass_0_in;
  wire PE_wrapper250_U0_fifo_cin_out_V_V_write_pass_0_out;
  wire [31:0] PE_wrapper250_U0_fifo_cout_drain_out_V_din_pass_0_out;
  wire fifo_cout_drain_PE_8_4_V_full_n_pass_0_in;
  wire PE_wrapper250_U0_fifo_cout_drain_out_V_write_pass_0_out;
  wire [255:0] PE_wrapper298_U0_fifo_cin_out_V_V_din_pass_0_out;
  wire fifo_cin_PE_13_4_V_V_full_n_pass_0_in;
  wire PE_wrapper298_U0_fifo_cin_out_V_V_write_pass_0_out;
  wire [63:0] cout_drain_IO_L1_out_wrapper432_U0_fifo_cout_drain_out_V_V_din_pass_0_in;
  wire fifo_cout_drain_cout_drain_IO_L1_out_4_14_V_V_full_n_pass_0_out;
  wire cout_drain_IO_L1_out_wrapper432_U0_fifo_cout_drain_out_V_V_write_pass_0_in;
  wire [255:0] PE_wrapper318_U0_fifo_w_out_V_V_din_pass_0_in;
  wire fifo_w_PE_14_1_V_V_full_n_pass_0_out;
  wire PE_wrapper318_U0_fifo_w_out_V_V_write_pass_0_in;
  wire [31:0] PE_wrapper306_U0_fifo_cout_drain_out_V_din_pass_0_in;
  wire fifo_cout_drain_PE_13_0_V_full_n_pass_0_out;
  wire PE_wrapper306_U0_fifo_cout_drain_out_V_write_pass_0_in;
  wire [31:0] PE_wrapper310_U0_fifo_cout_drain_out_V_din_pass_1_in;
  wire fifo_cout_drain_PE_13_4_V_full_n_pass_1_out;
  wire PE_wrapper310_U0_fifo_cout_drain_out_V_write_pass_1_in;
  wire [255:0] PE_wrapper286_U0_fifo_cin_out_V_V_din_pass_0_in;
  wire fifo_cin_PE_12_4_V_V_full_n_pass_0_out;
  wire PE_wrapper286_U0_fifo_cin_out_V_V_write_pass_0_in;
  wire [255:0] PE_wrapper331_U0_fifo_w_out_V_V_din_pass_0_out;
  wire fifo_w_PE_15_2_V_V_full_n_pass_0_in;
  wire PE_wrapper331_U0_fifo_w_out_V_V_write_pass_0_out;
  wire [31:0] PE_wrapper308_U0_fifo_cout_drain_out_V_din_pass_1_in;
  wire fifo_cout_drain_PE_13_2_V_full_n_pass_1_out;
  wire PE_wrapper308_U0_fifo_cout_drain_out_V_write_pass_1_in;
  wire [255:0] PE_wrapper330_U0_fifo_w_out_V_V_din_pass_0_in;
  wire fifo_w_PE_15_1_V_V_full_n_pass_0_out;
  wire PE_wrapper330_U0_fifo_w_out_V_V_write_pass_0_in;
  wire [255:0] PE_wrapper330_U0_fifo_cin_out_V_V_din_pass_0_in;
  wire fifo_cin_PE_16_0_V_V_full_n_pass_0_out;
  wire PE_wrapper330_U0_fifo_cin_out_V_V_write_pass_0_in;
  wire [63:0] cout_drain_IO_L1_out_wrapper419_U0_fifo_cout_drain_out_V_V_din_pass_0_in;
  wire fifo_cout_drain_cout_drain_IO_L1_out_3_11_V_V_full_n_pass_0_out;
  wire cout_drain_IO_L1_out_wrapper419_U0_fifo_cout_drain_out_V_V_write_pass_0_in;
  wire [255:0] w_IO_L2_in_boundary_U0_fifo_w_local_out_V_V_din_pass_0_out;
  wire fifo_w_PE_15_0_V_V_full_n_pass_0_in;
  wire w_IO_L2_in_boundary_U0_fifo_w_local_out_V_V_write_pass_0_out;
  wire [31:0] PE_wrapper333_U0_fifo_cout_drain_out_V_din_pass_0_in;
  wire fifo_cout_drain_PE_15_3_V_full_n_pass_0_out;
  wire PE_wrapper333_U0_fifo_cout_drain_out_V_write_pass_0_in;
  wire [255:0] PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_1_in;
  wire fifo_cin_PE_8_4_V_V_full_n_pass_1_out;
  wire PE_wrapper238_U0_fifo_cin_out_V_V_write_pass_1_in;
  wire [255:0] PE_wrapper297_U0_fifo_w_out_V_V_din_pass_1_in;
  wire fifo_w_PE_12_4_V_V_full_n_pass_1_out;
  wire PE_wrapper297_U0_fifo_w_out_V_V_write_pass_1_in;
  wire [255:0] PE_wrapper273_U0_fifo_w_out_V_V_din_pass_0_out;
  wire fifo_w_PE_10_4_V_V_full_n_pass_0_in;
  wire PE_wrapper273_U0_fifo_w_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_1_in;
  wire fifo_cin_PE_14_4_V_V_full_n_pass_1_out;
  wire PE_wrapper310_U0_fifo_cin_out_V_V_write_pass_1_in;
  wire [63:0] cout_drain_IO_L1_out_boundary_wrapper383_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_1_15_V_V_full_n_pass_0_in;
  wire cout_drain_IO_L1_out_boundary_wrapper383_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_1_in;
  wire fifo_cin_PE_14_1_V_V_full_n_pass_1_out;
  wire PE_wrapper307_U0_fifo_cin_out_V_V_write_pass_1_in;
  wire [31:0] PE_wrapper330_U0_fifo_cout_drain_out_V_din_pass_0_in;
  wire fifo_cout_drain_PE_15_0_V_full_n_pass_0_out;
  wire PE_wrapper330_U0_fifo_cout_drain_out_V_write_pass_0_in;
  wire [255:0] PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0_out;
  wire fifo_w_PE_8_5_V_V_full_n_pass_0_in;
  wire PE_wrapper250_U0_fifo_w_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper273_U0_fifo_cin_out_V_V_din_pass_0_out;
  wire fifo_cin_PE_11_3_V_V_full_n_pass_0_in;
  wire PE_wrapper273_U0_fifo_cin_out_V_V_write_pass_0_out;
  wire [63:0] cout_drain_IO_L1_out_wrapper369_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_0_13_V_V_full_n_pass_0_in;
  wire cout_drain_IO_L1_out_wrapper369_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper319_U0_fifo_w_out_V_V_din_pass_0_out;
  wire fifo_w_PE_14_2_V_V_full_n_pass_0_in;
  wire PE_wrapper319_U0_fifo_w_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper249_U0_fifo_w_out_V_V_din_pass_1_in;
  wire fifo_w_PE_8_4_V_V_full_n_pass_1_out;
  wire PE_wrapper249_U0_fifo_w_out_V_V_write_pass_1_in;
  wire [31:0] PE_wrapper319_U0_fifo_cout_drain_out_V_din_pass_0_out;
  wire fifo_cout_drain_PE_14_1_V_full_n_pass_0_in;
  wire PE_wrapper319_U0_fifo_cout_drain_out_V_write_pass_0_out;
  wire [255:0] PE_wrapper298_U0_fifo_w_out_V_V_din_pass_0_out;
  wire fifo_w_PE_12_5_V_V_full_n_pass_0_in;
  wire PE_wrapper298_U0_fifo_w_out_V_V_write_pass_0_out;
  wire [31:0] PE_wrapper334_U0_fifo_cout_drain_out_V_din_pass_0_out;
  wire fifo_cout_drain_PE_15_4_V_full_n_pass_0_in;
  wire PE_wrapper334_U0_fifo_cout_drain_out_V_write_pass_0_out;
  wire [255:0] PE_wrapper322_U0_fifo_w_out_V_V_din_pass_0_out;
  wire fifo_w_PE_14_5_V_V_full_n_pass_0_in;
  wire PE_wrapper322_U0_fifo_w_out_V_V_write_pass_0_out;
  wire [63:0] cout_drain_IO_L1_out_boundary_wrapper415_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_3_15_V_V_full_n_pass_0_in;
  wire cout_drain_IO_L1_out_boundary_wrapper415_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  wire [63:0] cout_drain_IO_L1_out_wrapper420_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_3_10_V_V_full_n_pass_0_in;
  wire cout_drain_IO_L1_out_wrapper420_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  wire [31:0] PE_wrapper318_U0_fifo_cout_drain_out_V_din_pass_0_in;
  wire fifo_cout_drain_PE_14_0_V_full_n_pass_0_out;
  wire PE_wrapper318_U0_fifo_cout_drain_out_V_write_pass_0_in;
  wire [255:0] PE_wrapper321_U0_fifo_w_out_V_V_din_pass_0_in;
  wire fifo_w_PE_14_4_V_V_full_n_pass_0_out;
  wire PE_wrapper321_U0_fifo_w_out_V_V_write_pass_0_in;
  wire [31:0] PE_wrapper322_U0_fifo_cout_drain_out_V_din_pass_0_out;
  wire fifo_cout_drain_PE_14_4_V_full_n_pass_0_in;
  wire PE_wrapper322_U0_fifo_cout_drain_out_V_write_pass_0_out;
  wire [255:0] PE_wrapper334_U0_fifo_w_out_V_V_din_pass_0_out;
  wire fifo_w_PE_15_5_V_V_full_n_pass_0_in;
  wire PE_wrapper334_U0_fifo_w_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper272_U0_fifo_w_out_V_V_din_pass_1_in;
  wire fifo_w_PE_10_3_V_V_full_n_pass_1_out;
  wire PE_wrapper272_U0_fifo_w_out_V_V_write_pass_1_in;
  wire [255:0] PE_wrapper261_U0_fifo_cin_out_V_V_din_pass_1_in;
  wire fifo_cin_PE_10_3_V_V_full_n_pass_1_out;
  wire PE_wrapper261_U0_fifo_cin_out_V_V_write_pass_1_in;
  wire [63:0] cout_drain_IO_L1_out_boundary_wrapper399_U0_fifo_cout_drain_out_V_V_din_pass_0_in;
  wire fifo_cout_drain_cout_drain_IO_L1_out_2_15_V_V_full_n_pass_0_out;
  wire cout_drain_IO_L1_out_boundary_wrapper399_U0_fifo_cout_drain_out_V_V_write_pass_0_in;
  wire [63:0] cout_drain_IO_L1_out_wrapper401_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_2_13_V_V_full_n_pass_0_in;
  wire cout_drain_IO_L1_out_wrapper401_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  wire [31:0] PE_wrapper298_U0_fifo_cout_drain_out_V_din_pass_0_out;
  wire fifo_cout_drain_PE_12_4_V_full_n_pass_0_in;
  wire PE_wrapper298_U0_fifo_cout_drain_out_V_write_pass_0_out;
  wire ap_start_Boundary_X2Y4_To_X4Y4_in;
  wire ap_rst_n_Boundary_X2Y4_To_X4Y4_in;
  wire ap_done_Boundary_X2Y4_To_X4Y4_out;
  wire ap_start_Boundary_X2Y6_To_X4Y6_out;
  wire ap_rst_n_Boundary_X2Y6_To_X4Y6_out;
  wire ap_done_Boundary_X2Y6_To_X4Y6_in;
  wire [31:0] PE_wrapper310_U0_fifo_cout_drain_out_V_din_pass_0_in;
  wire [31:0] PE_wrapper310_U0_fifo_cout_drain_out_V_din_pass_1_out;
  wire fifo_cout_drain_PE_13_4_V_full_n_pass_0_out;
  wire fifo_cout_drain_PE_13_4_V_full_n_pass_1_in;
  wire PE_wrapper310_U0_fifo_cout_drain_out_V_write_pass_0_in;
  wire PE_wrapper310_U0_fifo_cout_drain_out_V_write_pass_1_out;
  wire [31:0] PE_wrapper308_U0_fifo_cout_drain_out_V_din_pass_0_in;
  wire [31:0] PE_wrapper308_U0_fifo_cout_drain_out_V_din_pass_1_out;
  wire fifo_cout_drain_PE_13_2_V_full_n_pass_0_out;
  wire fifo_cout_drain_PE_13_2_V_full_n_pass_1_in;
  wire PE_wrapper308_U0_fifo_cout_drain_out_V_write_pass_0_in;
  wire PE_wrapper308_U0_fifo_cout_drain_out_V_write_pass_1_out;
  wire [255:0] PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0_in;
  wire [255:0] PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_1_out;
  wire fifo_cin_PE_8_4_V_V_full_n_pass_0_out;
  wire fifo_cin_PE_8_4_V_V_full_n_pass_1_in;
  wire PE_wrapper238_U0_fifo_cin_out_V_V_write_pass_0_in;
  wire PE_wrapper238_U0_fifo_cin_out_V_V_write_pass_1_out;
  wire [255:0] PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0_in;
  wire [255:0] PE_wrapper297_U0_fifo_w_out_V_V_din_pass_1_out;
  wire fifo_w_PE_12_4_V_V_full_n_pass_0_out;
  wire fifo_w_PE_12_4_V_V_full_n_pass_1_in;
  wire PE_wrapper297_U0_fifo_w_out_V_V_write_pass_0_in;
  wire PE_wrapper297_U0_fifo_w_out_V_V_write_pass_1_out;
  wire [255:0] PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0_in;
  wire [255:0] PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_1_out;
  wire fifo_cin_PE_14_4_V_V_full_n_pass_0_out;
  wire fifo_cin_PE_14_4_V_V_full_n_pass_1_in;
  wire PE_wrapper310_U0_fifo_cin_out_V_V_write_pass_0_in;
  wire PE_wrapper310_U0_fifo_cin_out_V_V_write_pass_1_out;
  wire [255:0] PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0_in;
  wire [255:0] PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_1_out;
  wire fifo_cin_PE_14_1_V_V_full_n_pass_0_out;
  wire fifo_cin_PE_14_1_V_V_full_n_pass_1_in;
  wire PE_wrapper307_U0_fifo_cin_out_V_V_write_pass_0_in;
  wire PE_wrapper307_U0_fifo_cin_out_V_V_write_pass_1_out;
  wire [255:0] PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0_in;
  wire [255:0] PE_wrapper250_U0_fifo_w_out_V_V_din_pass_1_out;
  wire fifo_w_PE_8_5_V_V_full_n_pass_0_out;
  wire fifo_w_PE_8_5_V_V_full_n_pass_1_in;
  wire PE_wrapper250_U0_fifo_w_out_V_V_write_pass_0_in;
  wire PE_wrapper250_U0_fifo_w_out_V_V_write_pass_1_out;
  wire [255:0] PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0_in;
  wire [255:0] PE_wrapper238_U0_fifo_w_out_V_V_din_pass_1_out;
  wire fifo_w_PE_7_5_V_V_full_n_pass_0_out;
  wire fifo_w_PE_7_5_V_V_full_n_pass_1_in;
  wire PE_wrapper238_U0_fifo_w_out_V_V_write_pass_0_in;
  wire PE_wrapper238_U0_fifo_w_out_V_V_write_pass_1_out;
  wire [31:0] PE_wrapper320_U0_fifo_cout_drain_out_V_din_pass_0_out;
  wire fifo_cout_drain_PE_14_2_V_full_n_pass_0_in;
  wire PE_wrapper320_U0_fifo_cout_drain_out_V_write_pass_0_out;
  wire [63:0] cout_drain_IO_L1_out_wrapper433_U0_fifo_cout_drain_out_V_V_din_pass_0_in;
  wire fifo_cout_drain_cout_drain_IO_L1_out_4_13_V_V_full_n_pass_0_out;
  wire cout_drain_IO_L1_out_wrapper433_U0_fifo_cout_drain_out_V_V_write_pass_0_in;
  wire [255:0] PE_wrapper309_U0_fifo_cin_out_V_V_din_pass_1_in;
  wire fifo_cin_PE_14_3_V_V_full_n_pass_1_out;
  wire PE_wrapper309_U0_fifo_cin_out_V_V_write_pass_1_in;
  wire [63:0] cout_drain_IO_L1_out_wrapper402_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_2_12_V_V_full_n_pass_0_in;
  wire cout_drain_IO_L1_out_wrapper402_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  wire [255:0] w_IO_L2_in149_U0_fifo_w_out_V_V_din_pass_0_out;
  wire fifo_w_w_IO_L2_in_15_V_V_full_n_pass_0_in;
  wire w_IO_L2_in149_U0_fifo_w_out_V_V_write_pass_0_out;
  wire [31:0] PE_wrapper286_U0_fifo_cout_drain_out_V_din_pass_0_out;
  wire fifo_cout_drain_PE_11_4_V_full_n_pass_0_in;
  wire PE_wrapper286_U0_fifo_cout_drain_out_V_write_pass_0_out;
  wire [255:0] PE_wrapper214_U0_fifo_cin_out_V_V_din_pass_1_in;
  wire fifo_cin_PE_6_4_V_V_full_n_pass_1_out;
  wire PE_wrapper214_U0_fifo_cin_out_V_V_write_pass_1_in;
  wire [63:0] cout_drain_IO_L1_out_wrapper432_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_4_14_V_V_full_n_pass_0_in;
  wire cout_drain_IO_L1_out_wrapper432_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper318_U0_fifo_w_out_V_V_din_pass_0_out;
  wire fifo_w_PE_14_1_V_V_full_n_pass_0_in;
  wire PE_wrapper318_U0_fifo_w_out_V_V_write_pass_0_out;
  wire [31:0] PE_wrapper226_U0_fifo_cout_drain_out_V_din_pass_0_out;
  wire fifo_cout_drain_PE_6_4_V_full_n_pass_0_in;
  wire PE_wrapper226_U0_fifo_cout_drain_out_V_write_pass_0_out;
  wire [255:0] PE_wrapper286_U0_fifo_cin_out_V_V_din_pass_0_out;
  wire fifo_cin_PE_12_4_V_V_full_n_pass_0_in;
  wire PE_wrapper286_U0_fifo_cin_out_V_V_write_pass_0_out;
  wire [255:0] w_IO_L2_in148_U0_fifo_w_out_V_V_din_pass_0_in;
  wire fifo_w_w_IO_L2_in_14_V_V_full_n_pass_0_out;
  wire w_IO_L2_in148_U0_fifo_w_out_V_V_write_pass_0_in;
  wire [255:0] PE_wrapper320_U0_fifo_cin_out_V_V_din_pass_0_out;
  wire fifo_cin_PE_15_2_V_V_full_n_pass_0_in;
  wire PE_wrapper320_U0_fifo_cin_out_V_V_write_pass_0_out;
  wire [63:0] cout_drain_IO_L1_out_wrapper418_U0_fifo_cout_drain_out_V_V_din_pass_1_in;
  wire fifo_cout_drain_cout_drain_IO_L1_out_3_12_V_V_full_n_pass_1_out;
  wire cout_drain_IO_L1_out_wrapper418_U0_fifo_cout_drain_out_V_V_write_pass_1_in;
  wire [255:0] PE_wrapper225_U0_fifo_w_out_V_V_din_pass_1_in;
  wire fifo_w_PE_6_4_V_V_full_n_pass_1_out;
  wire PE_wrapper225_U0_fifo_w_out_V_V_write_pass_1_in;
  wire [63:0] cout_drain_IO_L1_out_wrapper416_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_3_14_V_V_full_n_pass_0_in;
  wire cout_drain_IO_L1_out_wrapper416_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper330_U0_fifo_cin_out_V_V_din_pass_0_out;
  wire fifo_cin_PE_16_0_V_V_full_n_pass_0_in;
  wire PE_wrapper330_U0_fifo_cin_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper330_U0_fifo_w_out_V_V_din_pass_0_out;
  wire fifo_w_PE_15_1_V_V_full_n_pass_0_in;
  wire PE_wrapper330_U0_fifo_w_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper285_U0_fifo_w_out_V_V_din_pass_1_in;
  wire fifo_w_PE_11_4_V_V_full_n_pass_1_out;
  wire PE_wrapper285_U0_fifo_w_out_V_V_write_pass_1_in;
  wire [63:0] cout_drain_IO_L1_out_wrapper419_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_3_11_V_V_full_n_pass_0_in;
  wire cout_drain_IO_L1_out_wrapper419_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  wire [255:0] w_IO_L2_in_boundary_U0_fifo_w_local_out_V_V_din_pass_0_in;
  wire fifo_w_PE_15_0_V_V_full_n_pass_0_out;
  wire w_IO_L2_in_boundary_U0_fifo_w_local_out_V_V_write_pass_0_in;
  wire [255:0] PE_wrapper273_U0_fifo_w_out_V_V_din_pass_0_in;
  wire fifo_w_PE_10_4_V_V_full_n_pass_0_out;
  wire PE_wrapper273_U0_fifo_w_out_V_V_write_pass_0_in;
  wire [255:0] PE_wrapper286_U0_fifo_w_out_V_V_din_pass_0_out;
  wire fifo_w_PE_11_5_V_V_full_n_pass_0_in;
  wire PE_wrapper286_U0_fifo_w_out_V_V_write_pass_0_out;
  wire [63:0] cout_drain_IO_L1_out_boundary_wrapper383_U0_fifo_cout_drain_out_V_V_din_pass_0_in;
  wire fifo_cout_drain_cout_drain_IO_L1_out_1_15_V_V_full_n_pass_0_out;
  wire cout_drain_IO_L1_out_boundary_wrapper383_U0_fifo_cout_drain_out_V_V_write_pass_0_in;
  wire [31:0] PE_wrapper330_U0_fifo_cout_drain_out_V_din_pass_0_out;
  wire fifo_cout_drain_PE_15_0_V_full_n_pass_0_in;
  wire PE_wrapper330_U0_fifo_cout_drain_out_V_write_pass_0_out;
  wire [255:0] PE_wrapper306_U0_fifo_cin_out_V_V_din_pass_1_in;
  wire fifo_cin_PE_14_0_V_V_full_n_pass_1_out;
  wire PE_wrapper306_U0_fifo_cin_out_V_V_write_pass_1_in;
  wire [255:0] PE_wrapper321_U0_fifo_cin_out_V_V_din_pass_0_out;
  wire fifo_cin_PE_15_3_V_V_full_n_pass_0_in;
  wire PE_wrapper321_U0_fifo_cin_out_V_V_write_pass_0_out;
  wire [31:0] PE_wrapper285_U0_fifo_cout_drain_out_V_din_pass_1_in;
  wire fifo_cout_drain_PE_11_3_V_full_n_pass_1_out;
  wire PE_wrapper285_U0_fifo_cout_drain_out_V_write_pass_1_in;
  wire [255:0] PE_wrapper319_U0_fifo_w_out_V_V_din_pass_0_in;
  wire fifo_w_PE_14_2_V_V_full_n_pass_0_out;
  wire PE_wrapper319_U0_fifo_w_out_V_V_write_pass_0_in;
  wire [255:0] PE_wrapper226_U0_fifo_w_out_V_V_din_pass_0_out;
  wire fifo_w_PE_6_5_V_V_full_n_pass_0_in;
  wire PE_wrapper226_U0_fifo_w_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper308_U0_fifo_cin_out_V_V_din_pass_0_in;
  wire fifo_cin_PE_14_2_V_V_full_n_pass_0_out;
  wire PE_wrapper308_U0_fifo_cin_out_V_V_write_pass_0_in;
  wire [63:0] cout_drain_IO_L1_out_wrapper384_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_1_14_V_V_full_n_pass_0_in;
  wire cout_drain_IO_L1_out_wrapper384_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  wire [31:0] PE_wrapper319_U0_fifo_cout_drain_out_V_din_pass_0_in;
  wire fifo_cout_drain_PE_14_1_V_full_n_pass_0_out;
  wire PE_wrapper319_U0_fifo_cout_drain_out_V_write_pass_0_in;
  wire [31:0] PE_wrapper334_U0_fifo_cout_drain_out_V_din_pass_0_in;
  wire fifo_cout_drain_PE_15_4_V_full_n_pass_0_out;
  wire PE_wrapper334_U0_fifo_cout_drain_out_V_write_pass_0_in;
  wire [63:0] cout_drain_IO_L1_out_boundary_wrapper415_U0_fifo_cout_drain_out_V_V_din_pass_0_in;
  wire fifo_cout_drain_cout_drain_IO_L1_out_3_15_V_V_full_n_pass_0_out;
  wire cout_drain_IO_L1_out_boundary_wrapper415_U0_fifo_cout_drain_out_V_V_write_pass_0_in;
  wire [255:0] PE_wrapper274_U0_fifo_w_out_V_V_din_pass_0_out;
  wire fifo_w_PE_10_5_V_V_full_n_pass_0_in;
  wire PE_wrapper274_U0_fifo_w_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper262_U0_fifo_cin_out_V_V_din_pass_1_in;
  wire fifo_cin_PE_10_4_V_V_full_n_pass_1_out;
  wire PE_wrapper262_U0_fifo_cin_out_V_V_write_pass_1_in;
  wire [255:0] PE_wrapper226_U0_fifo_cin_out_V_V_din_pass_0_out;
  wire fifo_cin_PE_7_4_V_V_full_n_pass_0_in;
  wire PE_wrapper226_U0_fifo_cin_out_V_V_write_pass_0_out;
  wire [31:0] PE_wrapper318_U0_fifo_cout_drain_out_V_din_pass_0_out;
  wire fifo_cout_drain_PE_14_0_V_full_n_pass_0_in;
  wire PE_wrapper318_U0_fifo_cout_drain_out_V_write_pass_0_out;
  wire [31:0] PE_wrapper274_U0_fifo_cout_drain_out_V_din_pass_0_out;
  wire fifo_cout_drain_PE_10_4_V_full_n_pass_0_in;
  wire PE_wrapper274_U0_fifo_cout_drain_out_V_write_pass_0_out;
  wire [31:0] PE_wrapper296_U0_fifo_cout_drain_out_V_din_pass_1_in;
  wire fifo_cout_drain_PE_12_2_V_full_n_pass_1_out;
  wire PE_wrapper296_U0_fifo_cout_drain_out_V_write_pass_1_in;
  wire [255:0] PE_wrapper321_U0_fifo_w_out_V_V_din_pass_0_out;
  wire fifo_w_PE_14_4_V_V_full_n_pass_0_in;
  wire PE_wrapper321_U0_fifo_w_out_V_V_write_pass_0_out;
  wire [31:0] PE_wrapper322_U0_fifo_cout_drain_out_V_din_pass_0_in;
  wire fifo_cout_drain_PE_14_4_V_full_n_pass_0_out;
  wire PE_wrapper322_U0_fifo_cout_drain_out_V_write_pass_0_in;
  wire [63:0] cout_drain_IO_L1_out_wrapper401_U0_fifo_cout_drain_out_V_V_din_pass_0_in;
  wire fifo_cout_drain_cout_drain_IO_L1_out_2_13_V_V_full_n_pass_0_out;
  wire cout_drain_IO_L1_out_wrapper401_U0_fifo_cout_drain_out_V_V_write_pass_0_in;
  wire [63:0] cout_drain_IO_L1_out_wrapper434_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_4_12_V_V_full_n_pass_0_in;
  wire cout_drain_IO_L1_out_wrapper434_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  wire [31:0] PE_wrapper298_U0_fifo_cout_drain_out_V_din_pass_0_in;
  wire fifo_cout_drain_PE_12_4_V_full_n_pass_0_out;
  wire PE_wrapper298_U0_fifo_cout_drain_out_V_write_pass_0_in;
  wire ap_start_Boundary_X2Y6_To_X4Y6_in;
  wire ap_rst_n_Boundary_X2Y6_To_X4Y6_in;
  wire ap_done_Boundary_X2Y6_To_X4Y6_out;
  wire ap_start_Boundary_X2Y8_To_X4Y8_out;
  wire ap_rst_n_Boundary_X2Y8_To_X4Y8_out;
  wire ap_done_Boundary_X2Y8_To_X4Y8_in;
  wire [255:0] PE_wrapper288_U0_fifo_cin_out_V_V_din_pass_0_in;
  wire [255:0] PE_wrapper288_U0_fifo_cin_out_V_V_din_pass_1_out;
  wire fifo_cin_PE_12_6_V_V_full_n_pass_0_out;
  wire fifo_cin_PE_12_6_V_V_full_n_pass_1_in;
  wire PE_wrapper288_U0_fifo_cin_out_V_V_write_pass_0_in;
  wire PE_wrapper288_U0_fifo_cin_out_V_V_write_pass_1_out;
  wire [255:0] PE_wrapper311_U0_fifo_w_out_V_V_din_pass_0_out;
  wire fifo_w_PE_13_6_V_V_full_n_pass_0_in;
  wire PE_wrapper311_U0_fifo_w_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper251_U0_fifo_cin_out_V_V_din_pass_0_in;
  wire fifo_cin_PE_9_5_V_V_full_n_pass_0_out;
  wire PE_wrapper251_U0_fifo_cin_out_V_V_write_pass_0_in;
  wire [255:0] PE_wrapper299_U0_fifo_w_out_V_V_din_pass_0_out;
  wire fifo_w_PE_12_6_V_V_full_n_pass_0_in;
  wire PE_wrapper299_U0_fifo_w_out_V_V_write_pass_0_out;
  wire [31:0] PE_wrapper263_U0_fifo_cout_drain_out_V_din_pass_0_out;
  wire fifo_cout_drain_PE_9_5_V_full_n_pass_0_in;
  wire PE_wrapper263_U0_fifo_cout_drain_out_V_write_pass_0_out;
  wire [255:0] PE_wrapper310_U0_fifo_w_out_V_V_din_pass_0_in;
  wire fifo_w_PE_13_5_V_V_full_n_pass_0_out;
  wire PE_wrapper310_U0_fifo_w_out_V_V_write_pass_0_in;
  wire [31:0] PE_wrapper336_U0_fifo_cout_drain_out_V_din_pass_0_out;
  wire fifo_cout_drain_PE_15_6_V_full_n_pass_0_in;
  wire PE_wrapper336_U0_fifo_cout_drain_out_V_write_pass_0_out;
  wire [255:0] PE_wrapper262_U0_fifo_w_out_V_V_din_pass_1_in;
  wire fifo_w_PE_9_5_V_V_full_n_pass_1_out;
  wire PE_wrapper262_U0_fifo_w_out_V_V_write_pass_1_in;
  wire [255:0] PE_wrapper337_U0_fifo_w_out_V_V_din_pass_0_out;
  wire fifo_w_PE_15_8_V_V_full_n_pass_0_in;
  wire PE_wrapper337_U0_fifo_w_out_V_V_write_pass_0_out;
  wire [63:0] cout_drain_IO_L1_out_wrapper450_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_5_12_V_V_full_n_pass_0_in;
  wire cout_drain_IO_L1_out_wrapper450_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper298_U0_fifo_w_out_V_V_din_pass_2_in;
  wire fifo_w_PE_12_5_V_V_full_n_pass_2_out;
  wire PE_wrapper298_U0_fifo_w_out_V_V_write_pass_2_in;
  wire [255:0] PE_wrapper322_U0_fifo_w_out_V_V_din_pass_2_in;
  wire fifo_w_PE_14_5_V_V_full_n_pass_2_out;
  wire PE_wrapper322_U0_fifo_w_out_V_V_write_pass_2_in;
  wire [255:0] PE_wrapper263_U0_fifo_w_out_V_V_din_pass_0_out;
  wire fifo_w_PE_9_6_V_V_full_n_pass_0_in;
  wire PE_wrapper263_U0_fifo_w_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper323_U0_fifo_w_out_V_V_din_pass_0_out;
  wire fifo_w_PE_14_6_V_V_full_n_pass_0_in;
  wire PE_wrapper323_U0_fifo_w_out_V_V_write_pass_0_out;
  wire [31:0] PE_wrapper337_U0_fifo_cout_drain_out_V_din_pass_0_out;
  wire fifo_cout_drain_PE_15_7_V_full_n_pass_0_in;
  wire PE_wrapper337_U0_fifo_cout_drain_out_V_write_pass_0_out;
  wire [255:0] PE_wrapper324_U0_fifo_cin_out_V_V_din_pass_0_in;
  wire fifo_cin_PE_15_6_V_V_full_n_pass_0_out;
  wire PE_wrapper324_U0_fifo_cin_out_V_V_write_pass_0_in;
  wire [255:0] PE_wrapper334_U0_fifo_w_out_V_V_din_pass_2_in;
  wire fifo_w_PE_15_5_V_V_full_n_pass_2_out;
  wire PE_wrapper334_U0_fifo_w_out_V_V_write_pass_2_in;
  wire [255:0] PE_wrapper263_U0_fifo_cin_out_V_V_din_pass_0_out;
  wire fifo_cin_PE_10_5_V_V_full_n_pass_0_in;
  wire PE_wrapper263_U0_fifo_cin_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper325_U0_fifo_cin_out_V_V_din_pass_0_in;
  wire fifo_cin_PE_15_7_V_V_full_n_pass_0_out;
  wire PE_wrapper325_U0_fifo_cin_out_V_V_write_pass_0_in;
  wire [255:0] PE_wrapper287_U0_fifo_cin_out_V_V_din_pass_0_in;
  wire fifo_cin_PE_12_5_V_V_full_n_pass_0_out;
  wire PE_wrapper287_U0_fifo_cin_out_V_V_write_pass_0_in;
  wire ap_start_Boundary_X0Y8_To_X2Y8_in;
  wire ap_rst_n_Boundary_X0Y8_To_X2Y8_in;
  wire ap_done_Boundary_X0Y8_To_X2Y8_out;
  wire ap_start_Boundary_X0Y10_To_X2Y10_out;
  wire ap_rst_n_Boundary_X0Y10_To_X2Y10_out;
  wire ap_done_Boundary_X0Y10_To_X2Y10_in;
  wire [255:0] PE_wrapper337_U0_fifo_w_out_V_V_din_pass_0_in;
  wire [255:0] PE_wrapper337_U0_fifo_w_out_V_V_din_pass_1_out;
  wire fifo_w_PE_15_8_V_V_full_n_pass_0_out;
  wire fifo_w_PE_15_8_V_V_full_n_pass_1_in;
  wire PE_wrapper337_U0_fifo_w_out_V_V_write_pass_0_in;
  wire PE_wrapper337_U0_fifo_w_out_V_V_write_pass_1_out;
  wire [255:0] PE_wrapper311_U0_fifo_w_out_V_V_din_pass_0_in;
  wire fifo_w_PE_13_6_V_V_full_n_pass_0_out;
  wire PE_wrapper311_U0_fifo_w_out_V_V_write_pass_0_in;
  wire [255:0] PE_wrapper299_U0_fifo_w_out_V_V_din_pass_0_in;
  wire fifo_w_PE_12_6_V_V_full_n_pass_0_out;
  wire PE_wrapper299_U0_fifo_w_out_V_V_write_pass_0_in;
  wire [255:0] PE_wrapper289_U0_fifo_cin_out_V_V_din_pass_0_in;
  wire fifo_cin_PE_12_7_V_V_full_n_pass_0_out;
  wire PE_wrapper289_U0_fifo_cin_out_V_V_write_pass_0_in;
  wire [63:0] cout_drain_IO_L1_out_wrapper466_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_6_12_V_V_full_n_pass_0_in;
  wire cout_drain_IO_L1_out_wrapper466_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper290_U0_fifo_cin_out_V_V_din_pass_0_in;
  wire fifo_cin_PE_12_8_V_V_full_n_pass_0_out;
  wire PE_wrapper290_U0_fifo_cin_out_V_V_write_pass_0_in;
  wire [255:0] PE_wrapper302_U0_fifo_w_out_V_V_din_pass_0_out;
  wire fifo_w_PE_12_9_V_V_full_n_pass_0_in;
  wire PE_wrapper302_U0_fifo_w_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper325_U0_fifo_w_out_V_V_din_pass_0_out;
  wire fifo_w_PE_14_8_V_V_full_n_pass_0_in;
  wire PE_wrapper325_U0_fifo_w_out_V_V_write_pass_0_out;
  wire [31:0] PE_wrapper336_U0_fifo_cout_drain_out_V_din_pass_0_in;
  wire fifo_cout_drain_PE_15_6_V_full_n_pass_0_out;
  wire PE_wrapper336_U0_fifo_cout_drain_out_V_write_pass_0_in;
  wire [31:0] PE_wrapper302_U0_fifo_cout_drain_out_V_din_pass_0_out;
  wire fifo_cout_drain_PE_12_8_V_full_n_pass_0_in;
  wire PE_wrapper302_U0_fifo_cout_drain_out_V_write_pass_0_out;
  wire [255:0] PE_wrapper302_U0_fifo_cin_out_V_V_din_pass_0_out;
  wire fifo_cin_PE_13_8_V_V_full_n_pass_0_in;
  wire PE_wrapper302_U0_fifo_cin_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper288_U0_fifo_cin_out_V_V_din_pass_1_in;
  wire fifo_cin_PE_12_6_V_V_full_n_pass_1_out;
  wire PE_wrapper288_U0_fifo_cin_out_V_V_write_pass_1_in;
  wire [255:0] PE_wrapper323_U0_fifo_w_out_V_V_din_pass_0_in;
  wire fifo_w_PE_14_6_V_V_full_n_pass_0_out;
  wire PE_wrapper323_U0_fifo_w_out_V_V_write_pass_0_in;
  wire [31:0] PE_wrapper337_U0_fifo_cout_drain_out_V_din_pass_0_in;
  wire fifo_cout_drain_PE_15_7_V_full_n_pass_0_out;
  wire PE_wrapper337_U0_fifo_cout_drain_out_V_write_pass_0_in;
  wire [255:0] PE_wrapper324_U0_fifo_cin_out_V_V_din_pass_0_out;
  wire fifo_cin_PE_15_6_V_V_full_n_pass_0_in;
  wire PE_wrapper324_U0_fifo_cin_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper313_U0_fifo_w_out_V_V_din_pass_0_out;
  wire fifo_w_PE_13_8_V_V_full_n_pass_0_in;
  wire PE_wrapper313_U0_fifo_w_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper325_U0_fifo_cin_out_V_V_din_pass_0_out;
  wire fifo_cin_PE_15_7_V_V_full_n_pass_0_in;
  wire PE_wrapper325_U0_fifo_cin_out_V_V_write_pass_0_out;
  wire [63:0] cout_drain_IO_L1_out_wrapper482_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_7_12_V_V_full_n_pass_0_in;
  wire cout_drain_IO_L1_out_wrapper482_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  wire ap_start_Boundary_X0Y10_To_X2Y10_in;
  wire ap_rst_n_Boundary_X0Y10_To_X2Y10_in;
  wire ap_done_Boundary_X0Y10_To_X2Y10_out;
  wire ap_start_Boundary_X0Y12_To_X2Y12_out;
  wire ap_rst_n_Boundary_X0Y12_To_X2Y12_out;
  wire ap_done_Boundary_X0Y12_To_X2Y12_in;
  wire [255:0] PE_wrapper263_U0_fifo_w_out_V_V_din_pass_0_in;
  wire [255:0] PE_wrapper263_U0_fifo_w_out_V_V_din_pass_1_out;
  wire fifo_w_PE_9_6_V_V_full_n_pass_0_out;
  wire fifo_w_PE_9_6_V_V_full_n_pass_1_in;
  wire PE_wrapper263_U0_fifo_w_out_V_V_write_pass_0_in;
  wire PE_wrapper263_U0_fifo_w_out_V_V_write_pass_1_out;
  wire [255:0] PE_wrapper251_U0_fifo_cin_out_V_V_din_pass_0_out;
  wire fifo_cin_PE_9_5_V_V_full_n_pass_0_in;
  wire PE_wrapper251_U0_fifo_cin_out_V_V_write_pass_0_out;
  wire [31:0] PE_wrapper263_U0_fifo_cout_drain_out_V_din_pass_0_in;
  wire fifo_cout_drain_PE_9_5_V_full_n_pass_0_out;
  wire PE_wrapper263_U0_fifo_cout_drain_out_V_write_pass_0_in;
  wire [255:0] PE_wrapper276_U0_fifo_w_out_V_V_din_pass_0_out;
  wire fifo_w_PE_10_7_V_V_full_n_pass_0_in;
  wire PE_wrapper276_U0_fifo_w_out_V_V_write_pass_0_out;
  wire [31:0] PE_wrapper264_U0_fifo_cout_drain_out_V_din_pass_0_in;
  wire fifo_cout_drain_PE_9_6_V_full_n_pass_0_out;
  wire PE_wrapper264_U0_fifo_cout_drain_out_V_write_pass_0_in;
  wire [63:0] cout_drain_IO_L1_out_wrapper466_U0_fifo_cout_drain_out_V_V_din_pass_1_in;
  wire fifo_cout_drain_cout_drain_IO_L1_out_6_12_V_V_full_n_pass_1_out;
  wire cout_drain_IO_L1_out_wrapper466_U0_fifo_cout_drain_out_V_V_write_pass_1_in;
  wire [255:0] PE_wrapper264_U0_fifo_cin_out_V_V_din_pass_0_in;
  wire fifo_cin_PE_10_6_V_V_full_n_pass_0_out;
  wire PE_wrapper264_U0_fifo_cin_out_V_V_write_pass_0_in;
  wire [255:0] PE_wrapper286_U0_fifo_w_out_V_V_din_pass_0_in;
  wire fifo_w_PE_11_5_V_V_full_n_pass_0_out;
  wire PE_wrapper286_U0_fifo_w_out_V_V_write_pass_0_in;
  wire [255:0] PE_wrapper215_U0_fifo_cin_out_V_V_din_pass_0_in;
  wire fifo_cin_PE_6_5_V_V_full_n_pass_0_out;
  wire PE_wrapper215_U0_fifo_cin_out_V_V_write_pass_0_in;
  wire [255:0] PE_wrapper227_U0_fifo_w_out_V_V_din_pass_0_out;
  wire fifo_w_PE_6_6_V_V_full_n_pass_0_in;
  wire PE_wrapper227_U0_fifo_w_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper250_U0_fifo_w_out_V_V_din_pass_1_in;
  wire fifo_w_PE_8_5_V_V_full_n_pass_1_out;
  wire PE_wrapper250_U0_fifo_w_out_V_V_write_pass_1_in;
  wire [63:0] cout_drain_IO_L1_out_wrapper450_U0_fifo_cout_drain_out_V_V_din_pass_0_in;
  wire fifo_cout_drain_cout_drain_IO_L1_out_5_12_V_V_full_n_pass_0_out;
  wire cout_drain_IO_L1_out_wrapper450_U0_fifo_cout_drain_out_V_V_write_pass_0_in;
  wire [255:0] PE_wrapper226_U0_fifo_w_out_V_V_din_pass_0_in;
  wire fifo_w_PE_6_5_V_V_full_n_pass_0_out;
  wire PE_wrapper226_U0_fifo_w_out_V_V_write_pass_0_in;
  wire [63:0] cout_drain_IO_L1_out_wrapper456_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_5_6_V_V_full_n_pass_0_in;
  wire cout_drain_IO_L1_out_wrapper456_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper288_U0_fifo_cin_out_V_V_din_pass_0_out;
  wire fifo_cin_PE_12_6_V_V_full_n_pass_0_in;
  wire PE_wrapper288_U0_fifo_cin_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper251_U0_fifo_w_out_V_V_din_pass_0_out;
  wire fifo_w_PE_8_6_V_V_full_n_pass_0_in;
  wire PE_wrapper251_U0_fifo_w_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper274_U0_fifo_w_out_V_V_din_pass_0_in;
  wire fifo_w_PE_10_5_V_V_full_n_pass_0_out;
  wire PE_wrapper274_U0_fifo_w_out_V_V_write_pass_0_in;
  wire [255:0] PE_wrapper239_U0_fifo_w_out_V_V_din_pass_0_out;
  wire fifo_w_PE_7_6_V_V_full_n_pass_0_in;
  wire PE_wrapper239_U0_fifo_w_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper238_U0_fifo_w_out_V_V_din_pass_1_in;
  wire fifo_w_PE_7_5_V_V_full_n_pass_1_out;
  wire PE_wrapper238_U0_fifo_w_out_V_V_write_pass_1_in;
  wire [255:0] PE_wrapper263_U0_fifo_cin_out_V_V_din_pass_0_in;
  wire fifo_cin_PE_10_5_V_V_full_n_pass_0_out;
  wire PE_wrapper263_U0_fifo_cin_out_V_V_write_pass_0_in;
  wire [63:0] cout_drain_IO_L1_out_wrapper469_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_6_9_V_V_full_n_pass_0_in;
  wire cout_drain_IO_L1_out_wrapper469_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper288_U0_fifo_w_out_V_V_din_pass_0_out;
  wire fifo_w_PE_11_7_V_V_full_n_pass_0_in;
  wire PE_wrapper288_U0_fifo_w_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper287_U0_fifo_cin_out_V_V_din_pass_0_out;
  wire fifo_cin_PE_12_5_V_V_full_n_pass_0_in;
  wire PE_wrapper287_U0_fifo_cin_out_V_V_write_pass_0_out;
  wire ap_start_Boundary_X2Y8_To_X4Y8_in;
  wire ap_rst_n_Boundary_X2Y8_To_X4Y8_in;
  wire ap_done_Boundary_X2Y8_To_X4Y8_out;
  wire ap_start_Boundary_X2Y10_To_X4Y10_out;
  wire ap_rst_n_Boundary_X2Y10_To_X4Y10_out;
  wire ap_done_Boundary_X2Y10_To_X4Y10_in;
  wire [63:0] cout_drain_IO_L1_out_wrapper466_U0_fifo_cout_drain_out_V_V_din_pass_0_in;
  wire [63:0] cout_drain_IO_L1_out_wrapper466_U0_fifo_cout_drain_out_V_V_din_pass_1_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_6_12_V_V_full_n_pass_0_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_6_12_V_V_full_n_pass_1_in;
  wire cout_drain_IO_L1_out_wrapper466_U0_fifo_cout_drain_out_V_V_write_pass_0_in;
  wire cout_drain_IO_L1_out_wrapper466_U0_fifo_cout_drain_out_V_V_write_pass_1_out;
  wire [255:0] PE_wrapper302_U0_fifo_w_out_V_V_din_pass_0_in;
  wire [255:0] PE_wrapper302_U0_fifo_w_out_V_V_din_pass_1_out;
  wire fifo_w_PE_12_9_V_V_full_n_pass_0_out;
  wire fifo_w_PE_12_9_V_V_full_n_pass_1_in;
  wire PE_wrapper302_U0_fifo_w_out_V_V_write_pass_0_in;
  wire PE_wrapper302_U0_fifo_w_out_V_V_write_pass_1_out;
  wire [255:0] PE_wrapper290_U0_fifo_w_out_V_V_din_pass_0_out;
  wire fifo_w_PE_11_9_V_V_full_n_pass_0_in;
  wire PE_wrapper290_U0_fifo_w_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper253_U0_fifo_cin_out_V_V_din_pass_0_in;
  wire fifo_cin_PE_9_7_V_V_full_n_pass_0_out;
  wire PE_wrapper253_U0_fifo_cin_out_V_V_write_pass_0_in;
  wire [255:0] PE_wrapper289_U0_fifo_cin_out_V_V_din_pass_0_out;
  wire fifo_cin_PE_12_7_V_V_full_n_pass_0_in;
  wire PE_wrapper289_U0_fifo_cin_out_V_V_write_pass_0_out;
  wire [63:0] cout_drain_IO_L1_out_wrapper482_U0_fifo_cout_drain_out_V_V_din_pass_0_in;
  wire fifo_cout_drain_cout_drain_IO_L1_out_7_12_V_V_full_n_pass_0_out;
  wire cout_drain_IO_L1_out_wrapper482_U0_fifo_cout_drain_out_V_V_write_pass_0_in;
  wire [255:0] PE_wrapper276_U0_fifo_w_out_V_V_din_pass_0_in;
  wire fifo_w_PE_10_7_V_V_full_n_pass_0_out;
  wire PE_wrapper276_U0_fifo_w_out_V_V_write_pass_0_in;
  wire [31:0] PE_wrapper264_U0_fifo_cout_drain_out_V_din_pass_0_out;
  wire fifo_cout_drain_PE_9_6_V_full_n_pass_0_in;
  wire PE_wrapper264_U0_fifo_cout_drain_out_V_write_pass_0_out;
  wire [255:0] PE_wrapper278_U0_fifo_w_out_V_V_din_pass_0_out;
  wire fifo_w_PE_10_9_V_V_full_n_pass_0_in;
  wire PE_wrapper278_U0_fifo_w_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper290_U0_fifo_cin_out_V_V_din_pass_0_out;
  wire fifo_cin_PE_12_8_V_V_full_n_pass_0_in;
  wire PE_wrapper290_U0_fifo_cin_out_V_V_write_pass_0_out;
  wire [63:0] cout_drain_IO_L1_out_wrapper497_U0_fifo_cout_drain_out_V_V_din_pass_1_in;
  wire fifo_cout_drain_cout_drain_IO_L1_out_8_13_V_V_full_n_pass_1_out;
  wire cout_drain_IO_L1_out_wrapper497_U0_fifo_cout_drain_out_V_V_write_pass_1_in;
  wire [255:0] PE_wrapper264_U0_fifo_cin_out_V_V_din_pass_0_out;
  wire fifo_cin_PE_10_6_V_V_full_n_pass_0_in;
  wire PE_wrapper264_U0_fifo_cin_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper252_U0_fifo_cin_out_V_V_din_pass_0_in;
  wire fifo_cin_PE_9_6_V_V_full_n_pass_0_out;
  wire PE_wrapper252_U0_fifo_cin_out_V_V_write_pass_0_in;
  wire [31:0] PE_wrapper302_U0_fifo_cout_drain_out_V_din_pass_0_in;
  wire fifo_cout_drain_PE_12_8_V_full_n_pass_0_out;
  wire PE_wrapper302_U0_fifo_cout_drain_out_V_write_pass_0_in;
  wire [255:0] PE_wrapper266_U0_fifo_w_out_V_V_din_pass_0_out;
  wire fifo_w_PE_9_9_V_V_full_n_pass_0_in;
  wire PE_wrapper266_U0_fifo_w_out_V_V_write_pass_0_out;
  wire [63:0] cout_drain_IO_L1_out_wrapper501_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_8_9_V_V_full_n_pass_0_in;
  wire cout_drain_IO_L1_out_wrapper501_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper263_U0_fifo_w_out_V_V_din_pass_1_in;
  wire fifo_w_PE_9_6_V_V_full_n_pass_1_out;
  wire PE_wrapper263_U0_fifo_w_out_V_V_write_pass_1_in;
  wire [63:0] cout_drain_IO_L1_out_wrapper485_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_7_9_V_V_full_n_pass_0_in;
  wire cout_drain_IO_L1_out_wrapper485_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper254_U0_fifo_cin_out_V_V_din_pass_0_in;
  wire fifo_cin_PE_9_8_V_V_full_n_pass_0_out;
  wire PE_wrapper254_U0_fifo_cin_out_V_V_write_pass_0_in;
  wire [255:0] PE_wrapper288_U0_fifo_w_out_V_V_din_pass_0_in;
  wire fifo_w_PE_11_7_V_V_full_n_pass_0_out;
  wire PE_wrapper288_U0_fifo_w_out_V_V_write_pass_0_in;
  wire ap_start_Boundary_X2Y10_To_X4Y10_in;
  wire ap_rst_n_Boundary_X2Y10_To_X4Y10_in;
  wire ap_done_Boundary_X2Y10_To_X4Y10_out;
  wire ap_start_Boundary_X2Y12_To_X4Y12_out;
  wire ap_rst_n_Boundary_X2Y12_To_X4Y12_out;
  wire ap_done_Boundary_X2Y12_To_X4Y12_in;
  wire [255:0] PE_wrapper304_U0_fifo_cin_out_V_V_din_pass_0_in;
  wire [255:0] PE_wrapper304_U0_fifo_cin_out_V_V_din_pass_1_out;
  wire fifo_cin_PE_13_10_V_V_full_n_pass_0_out;
  wire fifo_cin_PE_13_10_V_V_full_n_pass_1_in;
  wire PE_wrapper304_U0_fifo_cin_out_V_V_write_pass_0_in;
  wire PE_wrapper304_U0_fifo_cin_out_V_V_write_pass_1_out;
  wire [255:0] PE_wrapper305_U0_fifo_cin_out_V_V_din_pass_0_in;
  wire [255:0] PE_wrapper305_U0_fifo_cin_out_V_V_din_pass_1_out;
  wire fifo_cin_PE_13_11_V_V_full_n_pass_0_out;
  wire fifo_cin_PE_13_11_V_V_full_n_pass_1_in;
  wire PE_wrapper305_U0_fifo_cin_out_V_V_write_pass_0_in;
  wire PE_wrapper305_U0_fifo_cin_out_V_V_write_pass_1_out;
  wire [63:0] cout_drain_IO_L1_out_wrapper513_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_9_13_V_V_full_n_pass_0_in;
  wire cout_drain_IO_L1_out_wrapper513_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper303_U0_fifo_cin_out_V_V_din_pass_0_in;
  wire fifo_cin_PE_13_9_V_V_full_n_pass_0_out;
  wire PE_wrapper303_U0_fifo_cin_out_V_V_write_pass_0_in;
  wire [255:0] PE_wrapper327_U0_fifo_w_out_V_V_din_pass_0_out;
  wire fifo_w_PE_14_10_V_V_full_n_pass_0_in;
  wire PE_wrapper327_U0_fifo_w_out_V_V_write_pass_0_out;
  wire [63:0] cout_drain_IO_L1_out_wrapper497_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_8_13_V_V_full_n_pass_0_in;
  wire cout_drain_IO_L1_out_wrapper497_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper325_U0_fifo_w_out_V_V_din_pass_0_in;
  wire fifo_w_PE_14_8_V_V_full_n_pass_0_out;
  wire PE_wrapper325_U0_fifo_w_out_V_V_write_pass_0_in;
  wire [255:0] PE_wrapper315_U0_fifo_w_out_V_V_din_pass_0_out;
  wire fifo_w_PE_13_10_V_V_full_n_pass_0_in;
  wire PE_wrapper315_U0_fifo_w_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper302_U0_fifo_cin_out_V_V_din_pass_0_in;
  wire fifo_cin_PE_13_8_V_V_full_n_pass_0_out;
  wire PE_wrapper302_U0_fifo_cin_out_V_V_write_pass_0_in;
  wire [255:0] PE_wrapper337_U0_fifo_w_out_V_V_din_pass_1_in;
  wire fifo_w_PE_15_8_V_V_full_n_pass_1_out;
  wire PE_wrapper337_U0_fifo_w_out_V_V_write_pass_1_in;
  wire [255:0] PE_wrapper313_U0_fifo_w_out_V_V_din_pass_0_in;
  wire fifo_w_PE_13_8_V_V_full_n_pass_0_out;
  wire PE_wrapper313_U0_fifo_w_out_V_V_write_pass_0_in;
  wire [255:0] PE_wrapper339_U0_fifo_w_out_V_V_din_pass_0_out;
  wire fifo_w_PE_15_10_V_V_full_n_pass_0_in;
  wire PE_wrapper339_U0_fifo_w_out_V_V_write_pass_0_out;
  wire ap_start_Boundary_X0Y12_To_X2Y12_in;
  wire ap_rst_n_Boundary_X0Y12_To_X2Y12_in;
  wire ap_done_Boundary_X0Y12_To_X2Y12_out;
  wire ap_start_Boundary_X0Y14_To_X2Y14_out;
  wire ap_rst_n_Boundary_X0Y14_To_X2Y14_out;
  wire ap_done_Boundary_X0Y14_To_X2Y14_in;
  wire [255:0] PE_wrapper304_U0_fifo_cin_out_V_V_din_pass_1_in;
  wire fifo_cin_PE_13_10_V_V_full_n_pass_1_out;
  wire PE_wrapper304_U0_fifo_cin_out_V_V_write_pass_1_in;
  wire [255:0] PE_wrapper327_U0_fifo_w_out_V_V_din_pass_0_in;
  wire fifo_w_PE_14_10_V_V_full_n_pass_0_out;
  wire PE_wrapper327_U0_fifo_w_out_V_V_write_pass_0_in;
  wire [255:0] PE_wrapper315_U0_fifo_w_out_V_V_din_pass_0_in;
  wire fifo_w_PE_13_10_V_V_full_n_pass_0_out;
  wire PE_wrapper315_U0_fifo_w_out_V_V_write_pass_0_in;
  wire [63:0] cout_drain_IO_L1_out_wrapper529_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_10_13_V_V_full_n_pass_0_in;
  wire cout_drain_IO_L1_out_wrapper529_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper305_U0_fifo_cin_out_V_V_din_pass_1_in;
  wire fifo_cin_PE_13_11_V_V_full_n_pass_1_out;
  wire PE_wrapper305_U0_fifo_cin_out_V_V_write_pass_1_in;
  wire [255:0] PE_wrapper339_U0_fifo_w_out_V_V_din_pass_0_in;
  wire fifo_w_PE_15_10_V_V_full_n_pass_0_out;
  wire PE_wrapper339_U0_fifo_w_out_V_V_write_pass_0_in;
  wire [63:0] cout_drain_IO_L1_out_wrapper544_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_11_13_V_V_full_n_pass_0_in;
  wire cout_drain_IO_L1_out_wrapper544_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  wire ap_start_Boundary_X0Y14_To_X2Y14_in;
  wire ap_rst_n_Boundary_X0Y14_To_X2Y14_in;
  wire ap_done_Boundary_X0Y14_To_X2Y14_out;
  wire [63:0] cout_drain_IO_L1_out_wrapper497_U0_fifo_cout_drain_out_V_V_din_pass_0_in;
  wire [63:0] cout_drain_IO_L1_out_wrapper497_U0_fifo_cout_drain_out_V_V_din_pass_1_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_8_13_V_V_full_n_pass_0_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_8_13_V_V_full_n_pass_1_in;
  wire cout_drain_IO_L1_out_wrapper497_U0_fifo_cout_drain_out_V_V_write_pass_0_in;
  wire cout_drain_IO_L1_out_wrapper497_U0_fifo_cout_drain_out_V_V_write_pass_1_out;
  wire [255:0] PE_wrapper278_U0_fifo_w_out_V_V_din_pass_0_in;
  wire [255:0] PE_wrapper278_U0_fifo_w_out_V_V_din_pass_1_out;
  wire fifo_w_PE_10_9_V_V_full_n_pass_0_out;
  wire fifo_w_PE_10_9_V_V_full_n_pass_1_in;
  wire PE_wrapper278_U0_fifo_w_out_V_V_write_pass_0_in;
  wire PE_wrapper278_U0_fifo_w_out_V_V_write_pass_1_out;
  wire [255:0] PE_wrapper290_U0_fifo_w_out_V_V_din_pass_0_in;
  wire fifo_w_PE_11_9_V_V_full_n_pass_0_out;
  wire PE_wrapper290_U0_fifo_w_out_V_V_write_pass_0_in;
  wire [255:0] PE_wrapper304_U0_fifo_cin_out_V_V_din_pass_0_out;
  wire fifo_cin_PE_13_10_V_V_full_n_pass_0_in;
  wire PE_wrapper304_U0_fifo_cin_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper279_U0_fifo_cin_out_V_V_din_pass_0_in;
  wire fifo_cin_PE_11_9_V_V_full_n_pass_0_out;
  wire PE_wrapper279_U0_fifo_cin_out_V_V_write_pass_0_in;
  wire [255:0] PE_wrapper267_U0_fifo_cin_out_V_V_din_pass_0_out;
  wire fifo_cin_PE_10_9_V_V_full_n_pass_0_in;
  wire PE_wrapper267_U0_fifo_cin_out_V_V_write_pass_0_out;
  wire [31:0] PE_wrapper269_U0_fifo_cout_drain_out_V_din_pass_0_in;
  wire fifo_cout_drain_PE_9_11_V_full_n_pass_0_out;
  wire PE_wrapper269_U0_fifo_cout_drain_out_V_write_pass_0_in;
  wire [63:0] cout_drain_IO_L1_out_wrapper513_U0_fifo_cout_drain_out_V_V_din_pass_0_in;
  wire fifo_cout_drain_cout_drain_IO_L1_out_9_13_V_V_full_n_pass_0_out;
  wire cout_drain_IO_L1_out_wrapper513_U0_fifo_cout_drain_out_V_V_write_pass_0_in;
  wire [255:0] PE_wrapper292_U0_fifo_w_out_V_V_din_pass_0_in;
  wire fifo_w_PE_11_11_V_V_full_n_pass_0_out;
  wire PE_wrapper292_U0_fifo_w_out_V_V_write_pass_0_in;
  wire [31:0] PE_wrapper281_U0_fifo_cout_drain_out_V_din_pass_0_in;
  wire fifo_cout_drain_PE_10_11_V_full_n_pass_0_out;
  wire PE_wrapper281_U0_fifo_cout_drain_out_V_write_pass_0_in;
  wire [31:0] PE_wrapper280_U0_fifo_cout_drain_out_V_din_pass_0_in;
  wire fifo_cout_drain_PE_10_10_V_full_n_pass_0_out;
  wire PE_wrapper280_U0_fifo_cout_drain_out_V_write_pass_0_in;
  wire [255:0] PE_wrapper281_U0_fifo_cin_out_V_V_din_pass_0_in;
  wire fifo_cin_PE_11_11_V_V_full_n_pass_0_out;
  wire PE_wrapper281_U0_fifo_cin_out_V_V_write_pass_0_in;
  wire [255:0] PE_wrapper302_U0_fifo_w_out_V_V_din_pass_1_in;
  wire fifo_w_PE_12_9_V_V_full_n_pass_1_out;
  wire PE_wrapper302_U0_fifo_w_out_V_V_write_pass_1_in;
  wire [255:0] PE_wrapper291_U0_fifo_w_out_V_V_din_pass_0_out;
  wire fifo_w_PE_11_10_V_V_full_n_pass_0_in;
  wire PE_wrapper291_U0_fifo_w_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper255_U0_fifo_cin_out_V_V_din_pass_0_in;
  wire fifo_cin_PE_9_9_V_V_full_n_pass_0_out;
  wire PE_wrapper255_U0_fifo_cin_out_V_V_write_pass_0_in;
  wire [255:0] PE_wrapper292_U0_fifo_cin_out_V_V_din_pass_0_in;
  wire fifo_cin_PE_12_10_V_V_full_n_pass_0_out;
  wire PE_wrapper292_U0_fifo_cin_out_V_V_write_pass_0_in;
  wire [63:0] cout_drain_IO_L1_out_wrapper517_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_9_9_V_V_full_n_pass_0_in;
  wire cout_drain_IO_L1_out_wrapper517_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  wire [31:0] PE_wrapper268_U0_fifo_cout_drain_out_V_din_pass_0_in;
  wire fifo_cout_drain_PE_9_10_V_full_n_pass_0_out;
  wire PE_wrapper268_U0_fifo_cout_drain_out_V_write_pass_0_in;
  wire [255:0] PE_wrapper266_U0_fifo_w_out_V_V_din_pass_0_in;
  wire fifo_w_PE_9_9_V_V_full_n_pass_0_out;
  wire PE_wrapper266_U0_fifo_w_out_V_V_write_pass_0_in;
  wire [63:0] cout_drain_IO_L1_out_wrapper529_U0_fifo_cout_drain_out_V_V_din_pass_1_in;
  wire fifo_cout_drain_cout_drain_IO_L1_out_10_13_V_V_full_n_pass_1_out;
  wire cout_drain_IO_L1_out_wrapper529_U0_fifo_cout_drain_out_V_V_write_pass_1_in;
  wire [63:0] cout_drain_IO_L1_out_wrapper533_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_10_9_V_V_full_n_pass_0_in;
  wire cout_drain_IO_L1_out_wrapper533_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper267_U0_fifo_w_out_V_V_din_pass_0_out;
  wire fifo_w_PE_9_10_V_V_full_n_pass_0_in;
  wire PE_wrapper267_U0_fifo_w_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper305_U0_fifo_cin_out_V_V_din_pass_0_out;
  wire fifo_cin_PE_13_11_V_V_full_n_pass_0_in;
  wire PE_wrapper305_U0_fifo_cin_out_V_V_write_pass_0_out;
  wire [31:0] PE_wrapper292_U0_fifo_cout_drain_out_V_din_pass_0_in;
  wire fifo_cout_drain_PE_11_10_V_full_n_pass_0_out;
  wire PE_wrapper292_U0_fifo_cout_drain_out_V_write_pass_0_in;
  wire [63:0] cout_drain_IO_L1_out_wrapper548_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_11_9_V_V_full_n_pass_0_in;
  wire cout_drain_IO_L1_out_wrapper548_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  wire [31:0] PE_wrapper279_U0_fifo_cout_drain_out_V_din_pass_0_in;
  wire fifo_cout_drain_PE_10_9_V_full_n_pass_0_out;
  wire PE_wrapper279_U0_fifo_cout_drain_out_V_write_pass_0_in;
  wire [255:0] PE_wrapper303_U0_fifo_cin_out_V_V_din_pass_0_out;
  wire fifo_cin_PE_13_9_V_V_full_n_pass_0_in;
  wire PE_wrapper303_U0_fifo_cin_out_V_V_write_pass_0_out;
  wire [63:0] cout_drain_IO_L1_out_wrapper544_U0_fifo_cout_drain_out_V_V_din_pass_1_in;
  wire fifo_cout_drain_cout_drain_IO_L1_out_11_13_V_V_full_n_pass_1_out;
  wire cout_drain_IO_L1_out_wrapper544_U0_fifo_cout_drain_out_V_V_write_pass_1_in;
  wire ap_start_Boundary_X2Y12_To_X4Y12_in;
  wire ap_rst_n_Boundary_X2Y12_To_X4Y12_in;
  wire ap_done_Boundary_X2Y12_To_X4Y12_out;
  wire ap_start_Boundary_X2Y14_To_X4Y14_out;
  wire ap_rst_n_Boundary_X2Y14_To_X4Y14_out;
  wire ap_done_Boundary_X2Y14_To_X4Y14_in;
  wire [63:0] cout_drain_IO_L1_out_wrapper529_U0_fifo_cout_drain_out_V_V_din_pass_0_in;
  wire [63:0] cout_drain_IO_L1_out_wrapper529_U0_fifo_cout_drain_out_V_V_din_pass_1_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_10_13_V_V_full_n_pass_0_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_10_13_V_V_full_n_pass_1_in;
  wire cout_drain_IO_L1_out_wrapper529_U0_fifo_cout_drain_out_V_V_write_pass_0_in;
  wire cout_drain_IO_L1_out_wrapper529_U0_fifo_cout_drain_out_V_V_write_pass_1_out;
  wire [63:0] cout_drain_IO_L1_out_wrapper544_U0_fifo_cout_drain_out_V_V_din_pass_0_in;
  wire [63:0] cout_drain_IO_L1_out_wrapper544_U0_fifo_cout_drain_out_V_V_din_pass_1_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_11_13_V_V_full_n_pass_0_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_11_13_V_V_full_n_pass_1_in;
  wire cout_drain_IO_L1_out_wrapper544_U0_fifo_cout_drain_out_V_V_write_pass_0_in;
  wire cout_drain_IO_L1_out_wrapper544_U0_fifo_cout_drain_out_V_V_write_pass_1_out;
  wire [255:0] PE_wrapper279_U0_fifo_cin_out_V_V_din_pass_0_out;
  wire fifo_cin_PE_11_9_V_V_full_n_pass_0_in;
  wire PE_wrapper279_U0_fifo_cin_out_V_V_write_pass_0_out;
  wire [31:0] PE_wrapper269_U0_fifo_cout_drain_out_V_din_pass_0_out;
  wire fifo_cout_drain_PE_9_11_V_full_n_pass_0_in;
  wire PE_wrapper269_U0_fifo_cout_drain_out_V_write_pass_0_out;
  wire [255:0] PE_wrapper267_U0_fifo_cin_out_V_V_din_pass_0_in;
  wire fifo_cin_PE_10_9_V_V_full_n_pass_0_out;
  wire PE_wrapper267_U0_fifo_cin_out_V_V_write_pass_0_in;
  wire [255:0] PE_wrapper292_U0_fifo_w_out_V_V_din_pass_0_out;
  wire fifo_w_PE_11_11_V_V_full_n_pass_0_in;
  wire PE_wrapper292_U0_fifo_w_out_V_V_write_pass_0_out;
  wire [31:0] PE_wrapper281_U0_fifo_cout_drain_out_V_din_pass_0_out;
  wire fifo_cout_drain_PE_10_11_V_full_n_pass_0_in;
  wire PE_wrapper281_U0_fifo_cout_drain_out_V_write_pass_0_out;
  wire [31:0] PE_wrapper280_U0_fifo_cout_drain_out_V_din_pass_0_out;
  wire fifo_cout_drain_PE_10_10_V_full_n_pass_0_in;
  wire PE_wrapper280_U0_fifo_cout_drain_out_V_write_pass_0_out;
  wire [255:0] PE_wrapper278_U0_fifo_w_out_V_V_din_pass_1_in;
  wire fifo_w_PE_10_9_V_V_full_n_pass_1_out;
  wire PE_wrapper278_U0_fifo_w_out_V_V_write_pass_1_in;
  wire [255:0] PE_wrapper281_U0_fifo_cin_out_V_V_din_pass_0_out;
  wire fifo_cin_PE_11_11_V_V_full_n_pass_0_in;
  wire PE_wrapper281_U0_fifo_cin_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper256_U0_fifo_cin_out_V_V_din_pass_1_in;
  wire fifo_cin_PE_9_10_V_V_full_n_pass_1_out;
  wire PE_wrapper256_U0_fifo_cin_out_V_V_write_pass_1_in;
  wire [255:0] PE_wrapper291_U0_fifo_w_out_V_V_din_pass_0_in;
  wire fifo_w_PE_11_10_V_V_full_n_pass_0_out;
  wire PE_wrapper291_U0_fifo_w_out_V_V_write_pass_0_in;
  wire [255:0] PE_wrapper292_U0_fifo_cin_out_V_V_din_pass_0_out;
  wire fifo_cin_PE_12_10_V_V_full_n_pass_0_in;
  wire PE_wrapper292_U0_fifo_cin_out_V_V_write_pass_0_out;
  wire [31:0] PE_wrapper268_U0_fifo_cout_drain_out_V_din_pass_0_out;
  wire fifo_cout_drain_PE_9_10_V_full_n_pass_0_in;
  wire PE_wrapper268_U0_fifo_cout_drain_out_V_write_pass_0_out;
  wire [255:0] PE_wrapper257_U0_fifo_cin_out_V_V_din_pass_1_in;
  wire fifo_cin_PE_9_11_V_V_full_n_pass_1_out;
  wire PE_wrapper257_U0_fifo_cin_out_V_V_write_pass_1_in;
  wire [255:0] PE_wrapper267_U0_fifo_w_out_V_V_din_pass_0_in;
  wire fifo_w_PE_9_10_V_V_full_n_pass_0_out;
  wire PE_wrapper267_U0_fifo_w_out_V_V_write_pass_0_in;
  wire [31:0] PE_wrapper292_U0_fifo_cout_drain_out_V_din_pass_0_out;
  wire fifo_cout_drain_PE_11_10_V_full_n_pass_0_in;
  wire PE_wrapper292_U0_fifo_cout_drain_out_V_write_pass_0_out;
  wire [31:0] PE_wrapper279_U0_fifo_cout_drain_out_V_din_pass_0_out;
  wire fifo_cout_drain_PE_10_9_V_full_n_pass_0_in;
  wire PE_wrapper279_U0_fifo_cout_drain_out_V_write_pass_0_out;
  wire ap_start_Boundary_X2Y14_To_X4Y14_in;
  wire ap_rst_n_Boundary_X2Y14_To_X4Y14_in;
  wire ap_done_Boundary_X2Y14_To_X4Y14_out;
  wire [255:0] w_IO_L2_in140_U0_fifo_w_out_V_V_din_pass_0_in;
  wire [255:0] w_IO_L2_in140_U0_fifo_w_out_V_V_din_pass_1_out;
  wire fifo_w_w_IO_L2_in_6_V_V_full_n_pass_0_out;
  wire fifo_w_w_IO_L2_in_6_V_V_full_n_pass_1_in;
  wire w_IO_L2_in140_U0_fifo_w_out_V_V_write_pass_0_in;
  wire w_IO_L2_in140_U0_fifo_w_out_V_V_write_pass_1_out;
  wire [255:0] PE_wrapper210_U0_fifo_cin_out_V_V_din_pass_0_in;
  wire [255:0] PE_wrapper210_U0_fifo_cin_out_V_V_din_pass_1_out;
  wire fifo_cin_PE_6_0_V_V_full_n_pass_0_out;
  wire fifo_cin_PE_6_0_V_V_full_n_pass_1_in;
  wire PE_wrapper210_U0_fifo_cin_out_V_V_write_pass_0_in;
  wire PE_wrapper210_U0_fifo_cin_out_V_V_write_pass_1_out;
  wire [255:0] w_IO_L2_in138_U0_fifo_w_local_out_V_V_din_pass_0_in;
  wire [255:0] w_IO_L2_in138_U0_fifo_w_local_out_V_V_din_pass_1_out;
  wire fifo_w_PE_3_0_V_V_full_n_pass_0_out;
  wire fifo_w_PE_3_0_V_V_full_n_pass_1_in;
  wire w_IO_L2_in138_U0_fifo_w_local_out_V_V_write_pass_0_in;
  wire w_IO_L2_in138_U0_fifo_w_local_out_V_V_write_pass_1_out;
  wire [63:0] cout_drain_IO_L1_out_wrapper378_U0_fifo_cout_drain_out_V_V_din_pass_0_in;
  wire [63:0] cout_drain_IO_L1_out_wrapper378_U0_fifo_cout_drain_out_V_V_din_pass_1_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_0_4_V_V_full_n_pass_0_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_0_4_V_V_full_n_pass_1_in;
  wire cout_drain_IO_L1_out_wrapper378_U0_fifo_cout_drain_out_V_V_write_pass_0_in;
  wire cout_drain_IO_L1_out_wrapper378_U0_fifo_cout_drain_out_V_V_write_pass_1_out;
  wire [255:0] PE_wrapper201_U0_fifo_w_out_V_V_din_pass_0_in;
  wire [255:0] PE_wrapper201_U0_fifo_w_out_V_V_din_pass_1_out;
  wire fifo_w_PE_4_4_V_V_full_n_pass_0_out;
  wire fifo_w_PE_4_4_V_V_full_n_pass_1_in;
  wire PE_wrapper201_U0_fifo_w_out_V_V_write_pass_0_in;
  wire PE_wrapper201_U0_fifo_w_out_V_V_write_pass_1_out;
  wire [255:0] PE_wrapper213_U0_fifo_w_out_V_V_din_pass_1_in;
  wire [255:0] PE_wrapper213_U0_fifo_w_out_V_V_din_pass_2_out;
  wire fifo_w_PE_5_4_V_V_full_n_pass_1_out;
  wire fifo_w_PE_5_4_V_V_full_n_pass_2_in;
  wire PE_wrapper213_U0_fifo_w_out_V_V_write_pass_1_in;
  wire PE_wrapper213_U0_fifo_w_out_V_V_write_pass_2_out;
  wire [63:0] kernel0_entry12_U0_w_V_out_din_pass_0_in;
  wire [63:0] kernel0_entry12_U0_w_V_out_din_pass_1_out;
  wire w_V_c_full_n_pass_0_out;
  wire w_V_c_full_n_pass_1_in;
  wire kernel0_entry12_U0_w_V_out_write_pass_0_in;
  wire kernel0_entry12_U0_w_V_out_write_pass_1_out;
  wire [63:0] kernel0_entry12_U0_cout_V_out_din_pass_0_in;
  wire [63:0] kernel0_entry12_U0_cout_V_out_din_pass_1_out;
  wire cout_V_c_full_n_pass_0_out;
  wire cout_V_c_full_n_pass_1_in;
  wire kernel0_entry12_U0_cout_V_out_write_pass_0_in;
  wire kernel0_entry12_U0_cout_V_out_write_pass_1_out;
  wire [255:0] PE_wrapper165_U0_fifo_w_out_V_V_din_pass_0_out;
  wire fifo_w_PE_1_4_V_V_full_n_pass_0_in;
  wire PE_wrapper165_U0_fifo_w_out_V_V_write_pass_0_out;
  wire [255:0] cin_IO_L2_in127_U0_fifo_cin_out_V_V_din_pass_0_out;
  wire fifo_cin_cin_IO_L2_in_4_V_V_full_n_pass_0_in;
  wire cin_IO_L2_in127_U0_fifo_cin_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper163_U0_fifo_w_out_V_V_din_pass_0_in;
  wire fifo_w_PE_1_2_V_V_full_n_pass_0_out;
  wire PE_wrapper163_U0_fifo_w_out_V_V_write_pass_0_in;
  wire [255:0] PE_wrapper188_U0_fifo_w_out_V_V_din_pass_0_in;
  wire fifo_w_PE_3_3_V_V_full_n_pass_0_out;
  wire PE_wrapper188_U0_fifo_w_out_V_V_write_pass_0_in;
  wire [255:0] w_IO_L2_in136_U0_fifo_w_out_V_V_din_pass_0_out;
  wire fifo_w_w_IO_L2_in_2_V_V_full_n_pass_0_in;
  wire w_IO_L2_in136_U0_fifo_w_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper153_U0_fifo_w_out_V_V_din_pass_0_out;
  wire fifo_w_PE_0_4_V_V_full_n_pass_0_in;
  wire PE_wrapper153_U0_fifo_w_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper177_U0_fifo_w_out_V_V_din_pass_0_out;
  wire fifo_w_PE_2_4_V_V_full_n_pass_0_in;
  wire PE_wrapper177_U0_fifo_w_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper151_U0_fifo_w_out_V_V_din_pass_0_in;
  wire fifo_w_PE_0_2_V_V_full_n_pass_0_out;
  wire PE_wrapper151_U0_fifo_w_out_V_V_write_pass_0_in;
  wire [31:0] PE_wrapper165_U0_fifo_cout_drain_out_V_din_pass_0_out;
  wire fifo_cout_drain_PE_1_3_V_full_n_pass_0_in;
  wire PE_wrapper165_U0_fifo_cout_drain_out_V_write_pass_0_out;
  wire [255:0] PE_wrapper150_U0_fifo_cin_out_V_V_din_pass_0_in;
  wire fifo_cin_PE_1_0_V_V_full_n_pass_0_out;
  wire PE_wrapper150_U0_fifo_cin_out_V_V_write_pass_0_in;
  wire [31:0] PE_wrapper153_U0_fifo_cout_drain_out_V_din_pass_0_out;
  wire fifo_cout_drain_PE_0_3_V_full_n_pass_0_in;
  wire PE_wrapper153_U0_fifo_cout_drain_out_V_write_pass_0_out;
  wire [31:0] PE_wrapper177_U0_fifo_cout_drain_out_V_din_pass_0_out;
  wire fifo_cout_drain_PE_2_3_V_full_n_pass_0_in;
  wire PE_wrapper177_U0_fifo_cout_drain_out_V_write_pass_0_out;
  wire [31:0] PE_wrapper164_U0_fifo_cout_drain_out_V_din_pass_0_out;
  wire fifo_cout_drain_PE_1_2_V_full_n_pass_0_in;
  wire PE_wrapper164_U0_fifo_cout_drain_out_V_write_pass_0_out;
  wire [31:0] PE_wrapper189_U0_fifo_cout_drain_out_V_din_pass_0_out;
  wire fifo_cout_drain_PE_3_3_V_full_n_pass_0_in;
  wire PE_wrapper189_U0_fifo_cout_drain_out_V_write_pass_0_out;
  wire [255:0] PE_wrapper162_U0_fifo_cin_out_V_V_din_pass_0_out;
  wire fifo_cin_PE_2_0_V_V_full_n_pass_0_in;
  wire PE_wrapper162_U0_fifo_cin_out_V_V_write_pass_0_out;
  wire [255:0] w_IO_L3_in_serialize_U0_fifo_w_local_out_V_V_din_pass_0_in;
  wire fifo_w_w_IO_L3_in_serialize_V_V_full_n_pass_0_out;
  wire w_IO_L3_in_serialize_U0_fifo_w_local_out_V_V_write_pass_0_in;
  wire [255:0] cin_IO_L2_in125_U0_fifo_cin_out_V_V_din_pass_1_in;
  wire fifo_cin_cin_IO_L2_in_2_V_V_full_n_pass_1_out;
  wire cin_IO_L2_in125_U0_fifo_cin_out_V_V_write_pass_1_in;
  wire [31:0] PE_wrapper152_U0_fifo_cout_drain_out_V_din_pass_0_out;
  wire fifo_cout_drain_PE_0_2_V_full_n_pass_0_in;
  wire PE_wrapper152_U0_fifo_cout_drain_out_V_write_pass_0_out;
  wire [255:0] PE_wrapper189_U0_fifo_w_out_V_V_din_pass_0_out;
  wire fifo_w_PE_3_4_V_V_full_n_pass_0_in;
  wire PE_wrapper189_U0_fifo_w_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper175_U0_fifo_w_out_V_V_din_pass_0_in;
  wire fifo_w_PE_2_2_V_V_full_n_pass_0_out;
  wire PE_wrapper175_U0_fifo_w_out_V_V_write_pass_0_in;
  wire [255:0] PE_wrapper162_U0_fifo_w_out_V_V_din_pass_0_out;
  wire fifo_w_PE_1_1_V_V_full_n_pass_0_in;
  wire PE_wrapper162_U0_fifo_w_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper189_U0_fifo_cin_out_V_V_din_pass_0_out;
  wire fifo_cin_PE_4_3_V_V_full_n_pass_0_in;
  wire PE_wrapper189_U0_fifo_cin_out_V_V_write_pass_0_out;
  wire [31:0] PE_wrapper176_U0_fifo_cout_drain_out_V_din_pass_0_out;
  wire fifo_cout_drain_PE_2_2_V_full_n_pass_0_in;
  wire PE_wrapper176_U0_fifo_cout_drain_out_V_write_pass_0_out;
  wire [255:0] PE_wrapper176_U0_fifo_cin_out_V_V_din_pass_0_out;
  wire fifo_cin_PE_3_2_V_V_full_n_pass_0_in;
  wire PE_wrapper176_U0_fifo_cin_out_V_V_write_pass_0_out;
  wire [31:0] PE_wrapper162_U0_fifo_cout_drain_out_V_din_pass_0_out;
  wire fifo_cout_drain_PE_1_0_V_full_n_pass_0_in;
  wire PE_wrapper162_U0_fifo_cout_drain_out_V_write_pass_0_out;
  wire [255:0] w_IO_L2_in135_U0_fifo_w_local_out_V_V_din_pass_0_out;
  wire fifo_w_PE_0_0_V_V_full_n_pass_0_in;
  wire w_IO_L2_in135_U0_fifo_w_local_out_V_V_write_pass_0_out;
  wire ap_start_Boundary_X4Y2_To_X6Y2_in;
  wire ap_rst_n_Boundary_X4Y2_To_X6Y2_in;
  wire ap_done_Boundary_X4Y2_To_X6Y2_out;
  wire ap_start_Boundary_X4Y4_To_X6Y4_out;
  wire ap_rst_n_Boundary_X4Y4_To_X6Y4_out;
  wire ap_done_Boundary_X4Y4_To_X6Y4_in;
  wire [255:0] PE_wrapper187_U0_fifo_w_out_V_V_din_pass_0_in;
  wire [255:0] PE_wrapper187_U0_fifo_w_out_V_V_din_pass_1_out;
  wire fifo_w_PE_3_2_V_V_full_n_pass_0_out;
  wire fifo_w_PE_3_2_V_V_full_n_pass_1_in;
  wire PE_wrapper187_U0_fifo_w_out_V_V_write_pass_0_in;
  wire PE_wrapper187_U0_fifo_w_out_V_V_write_pass_1_out;
  wire [31:0] PE_wrapper163_U0_fifo_cout_drain_out_V_din_pass_0_in;
  wire [31:0] PE_wrapper163_U0_fifo_cout_drain_out_V_din_pass_1_out;
  wire fifo_cout_drain_PE_1_1_V_full_n_pass_0_out;
  wire fifo_cout_drain_PE_1_1_V_full_n_pass_1_in;
  wire PE_wrapper163_U0_fifo_cout_drain_out_V_write_pass_0_in;
  wire PE_wrapper163_U0_fifo_cout_drain_out_V_write_pass_1_out;
  wire [31:0] PE_wrapper175_U0_fifo_cout_drain_out_V_din_pass_0_in;
  wire [31:0] PE_wrapper175_U0_fifo_cout_drain_out_V_din_pass_1_out;
  wire fifo_cout_drain_PE_2_1_V_full_n_pass_0_out;
  wire fifo_cout_drain_PE_2_1_V_full_n_pass_1_in;
  wire PE_wrapper175_U0_fifo_cout_drain_out_V_write_pass_0_in;
  wire PE_wrapper175_U0_fifo_cout_drain_out_V_write_pass_1_out;
  wire [255:0] PE_wrapper187_U0_fifo_cin_out_V_V_din_pass_0_in;
  wire [255:0] PE_wrapper187_U0_fifo_cin_out_V_V_din_pass_1_out;
  wire fifo_cin_PE_4_1_V_V_full_n_pass_0_out;
  wire fifo_cin_PE_4_1_V_V_full_n_pass_1_in;
  wire PE_wrapper187_U0_fifo_cin_out_V_V_write_pass_0_in;
  wire PE_wrapper187_U0_fifo_cin_out_V_V_write_pass_1_out;
  wire [255:0] PE_wrapper186_U0_fifo_cin_out_V_V_din_pass_0_in;
  wire [255:0] PE_wrapper186_U0_fifo_cin_out_V_V_din_pass_1_out;
  wire fifo_cin_PE_4_0_V_V_full_n_pass_0_out;
  wire fifo_cin_PE_4_0_V_V_full_n_pass_1_in;
  wire PE_wrapper186_U0_fifo_cin_out_V_V_write_pass_0_in;
  wire PE_wrapper186_U0_fifo_cin_out_V_V_write_pass_1_out;
  wire [31:0] PE_wrapper187_U0_fifo_cout_drain_out_V_din_pass_0_in;
  wire [31:0] PE_wrapper187_U0_fifo_cout_drain_out_V_din_pass_1_out;
  wire fifo_cout_drain_PE_3_1_V_full_n_pass_0_out;
  wire fifo_cout_drain_PE_3_1_V_full_n_pass_1_in;
  wire PE_wrapper187_U0_fifo_cout_drain_out_V_write_pass_0_in;
  wire PE_wrapper187_U0_fifo_cout_drain_out_V_write_pass_1_out;
  wire [255:0] w_IO_L2_in137_U0_fifo_w_out_V_V_din_pass_0_in;
  wire [255:0] w_IO_L2_in137_U0_fifo_w_out_V_V_din_pass_1_out;
  wire fifo_w_w_IO_L2_in_3_V_V_full_n_pass_0_out;
  wire fifo_w_w_IO_L2_in_3_V_V_full_n_pass_1_in;
  wire w_IO_L2_in137_U0_fifo_w_out_V_V_write_pass_0_in;
  wire w_IO_L2_in137_U0_fifo_w_out_V_V_write_pass_1_out;
  wire [63:0] cout_drain_IO_L1_out_wrapper376_U0_fifo_cout_drain_out_V_V_din_pass_1_in;
  wire [63:0] cout_drain_IO_L1_out_wrapper376_U0_fifo_cout_drain_out_V_V_din_pass_2_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_0_6_V_V_full_n_pass_1_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_0_6_V_V_full_n_pass_2_in;
  wire cout_drain_IO_L1_out_wrapper376_U0_fifo_cout_drain_out_V_V_write_pass_1_in;
  wire cout_drain_IO_L1_out_wrapper376_U0_fifo_cout_drain_out_V_V_write_pass_2_out;
  wire [31:0] PE_wrapper151_U0_fifo_cout_drain_out_V_din_pass_0_in;
  wire [31:0] PE_wrapper151_U0_fifo_cout_drain_out_V_din_pass_1_out;
  wire fifo_cout_drain_PE_0_1_V_full_n_pass_0_out;
  wire fifo_cout_drain_PE_0_1_V_full_n_pass_1_in;
  wire PE_wrapper151_U0_fifo_cout_drain_out_V_write_pass_0_in;
  wire PE_wrapper151_U0_fifo_cout_drain_out_V_write_pass_1_out;
  wire [63:0] cout_drain_IO_L1_out_wrapper392_U0_fifo_cout_drain_out_V_V_din_pass_1_in;
  wire [63:0] cout_drain_IO_L1_out_wrapper392_U0_fifo_cout_drain_out_V_V_din_pass_2_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_1_6_V_V_full_n_pass_1_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_1_6_V_V_full_n_pass_2_in;
  wire cout_drain_IO_L1_out_wrapper392_U0_fifo_cout_drain_out_V_V_write_pass_1_in;
  wire cout_drain_IO_L1_out_wrapper392_U0_fifo_cout_drain_out_V_V_write_pass_2_out;
  wire [63:0] cout_drain_IO_L2_out564_U0_fifo_cout_drain_out_V_V_din_pass_1_in;
  wire fifo_cout_drain_cout_drain_IO_L2_out_4_V_V_full_n_pass_1_out;
  wire cout_drain_IO_L2_out564_U0_fifo_cout_drain_out_V_V_write_pass_1_in;
  wire [31:0] PE_wrapper200_U0_fifo_cout_drain_out_V_din_pass_0_in;
  wire fifo_cout_drain_PE_4_2_V_full_n_pass_0_out;
  wire PE_wrapper200_U0_fifo_cout_drain_out_V_write_pass_0_in;
  wire [255:0] PE_wrapper212_U0_fifo_cin_out_V_V_din_pass_0_out;
  wire fifo_cin_PE_6_2_V_V_full_n_pass_0_in;
  wire PE_wrapper212_U0_fifo_cin_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper210_U0_fifo_w_out_V_V_din_pass_0_in;
  wire fifo_w_PE_5_1_V_V_full_n_pass_0_out;
  wire PE_wrapper210_U0_fifo_w_out_V_V_write_pass_0_in;
  wire [31:0] PE_wrapper188_U0_fifo_cout_drain_out_V_din_pass_0_in;
  wire fifo_cout_drain_PE_3_2_V_full_n_pass_0_out;
  wire PE_wrapper188_U0_fifo_cout_drain_out_V_write_pass_0_in;
  wire [63:0] cout_drain_IO_L1_out_wrapper424_U0_fifo_cout_drain_out_V_V_din_pass_1_in;
  wire fifo_cout_drain_cout_drain_IO_L1_out_3_6_V_V_full_n_pass_1_out;
  wire cout_drain_IO_L1_out_wrapper424_U0_fifo_cout_drain_out_V_V_write_pass_1_in;
  wire [255:0] PE_wrapper201_U0_fifo_cin_out_V_V_din_pass_0_in;
  wire fifo_cin_PE_5_3_V_V_full_n_pass_0_out;
  wire PE_wrapper201_U0_fifo_cin_out_V_V_write_pass_0_in;
  wire [63:0] cout_drain_IO_L1_out_wrapper398_U0_fifo_cout_drain_out_V_V_din_pass_0_in;
  wire fifo_cout_drain_cout_drain_IO_L1_out_1_0_V_V_full_n_pass_0_out;
  wire cout_drain_IO_L1_out_wrapper398_U0_fifo_cout_drain_out_V_V_write_pass_0_in;
  wire [255:0] PE_wrapper199_U0_fifo_cin_out_V_V_din_pass_0_in;
  wire fifo_cin_PE_5_1_V_V_full_n_pass_0_out;
  wire PE_wrapper199_U0_fifo_cin_out_V_V_write_pass_0_in;
  wire [255:0] PE_wrapper211_U0_fifo_cin_out_V_V_din_pass_0_out;
  wire fifo_cin_PE_6_1_V_V_full_n_pass_0_in;
  wire PE_wrapper211_U0_fifo_cin_out_V_V_write_pass_0_out;
  wire [31:0] PE_wrapper165_U0_fifo_cout_drain_out_V_din_pass_1_in;
  wire fifo_cout_drain_PE_1_3_V_full_n_pass_1_out;
  wire PE_wrapper165_U0_fifo_cout_drain_out_V_write_pass_1_in;
  wire [31:0] PE_wrapper211_U0_fifo_cout_drain_out_V_din_pass_0_out;
  wire fifo_cout_drain_PE_5_1_V_full_n_pass_0_in;
  wire PE_wrapper211_U0_fifo_cout_drain_out_V_write_pass_0_out;
  wire [31:0] PE_wrapper153_U0_fifo_cout_drain_out_V_din_pass_1_in;
  wire fifo_cout_drain_PE_0_3_V_full_n_pass_1_out;
  wire PE_wrapper153_U0_fifo_cout_drain_out_V_write_pass_1_in;
  wire [31:0] PE_wrapper201_U0_fifo_cout_drain_out_V_din_pass_0_in;
  wire fifo_cout_drain_PE_4_3_V_full_n_pass_0_out;
  wire PE_wrapper201_U0_fifo_cout_drain_out_V_write_pass_0_in;
  wire [63:0] cout_drain_IO_L1_out_wrapper382_U0_fifo_cout_drain_out_V_V_din_pass_0_in;
  wire fifo_cout_drain_cout_drain_IO_L1_out_0_0_V_V_full_n_pass_0_out;
  wire cout_drain_IO_L1_out_wrapper382_U0_fifo_cout_drain_out_V_V_write_pass_0_in;
  wire [255:0] PE_wrapper213_U0_fifo_cin_out_V_V_din_pass_0_out;
  wire fifo_cin_PE_6_3_V_V_full_n_pass_0_in;
  wire PE_wrapper213_U0_fifo_cin_out_V_V_write_pass_0_out;
  wire [31:0] PE_wrapper177_U0_fifo_cout_drain_out_V_din_pass_1_in;
  wire fifo_cout_drain_PE_2_3_V_full_n_pass_1_out;
  wire PE_wrapper177_U0_fifo_cout_drain_out_V_write_pass_1_in;
  wire [31:0] PE_wrapper164_U0_fifo_cout_drain_out_V_din_pass_1_in;
  wire fifo_cout_drain_PE_1_2_V_full_n_pass_1_out;
  wire PE_wrapper164_U0_fifo_cout_drain_out_V_write_pass_1_in;
  wire [31:0] PE_wrapper189_U0_fifo_cout_drain_out_V_din_pass_1_in;
  wire fifo_cout_drain_PE_3_3_V_full_n_pass_1_out;
  wire PE_wrapper189_U0_fifo_cout_drain_out_V_write_pass_1_in;
  wire [255:0] cin_IO_L2_in124_U0_fifo_cin_out_V_V_din_pass_0_in;
  wire fifo_cin_cin_IO_L2_in_1_V_V_full_n_pass_0_out;
  wire cin_IO_L2_in124_U0_fifo_cin_out_V_V_write_pass_0_in;
  wire [31:0] PE_wrapper152_U0_fifo_cout_drain_out_V_din_pass_1_in;
  wire fifo_cout_drain_PE_0_2_V_full_n_pass_1_out;
  wire PE_wrapper152_U0_fifo_cout_drain_out_V_write_pass_1_in;
  wire [255:0] cin_IO_L2_in125_U0_fifo_cin_out_V_V_din_pass_0_out;
  wire fifo_cin_cin_IO_L2_in_2_V_V_full_n_pass_0_in;
  wire cin_IO_L2_in125_U0_fifo_cin_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper200_U0_fifo_cin_out_V_V_din_pass_0_in;
  wire fifo_cin_PE_5_2_V_V_full_n_pass_0_out;
  wire PE_wrapper200_U0_fifo_cin_out_V_V_write_pass_0_in;
  wire [255:0] cin_IO_L2_in125_U0_fifo_cin_local_out_V_V_din_pass_0_out;
  wire fifo_cin_PE_0_1_V_V_full_n_pass_0_in;
  wire cin_IO_L2_in125_U0_fifo_cin_local_out_V_V_write_pass_0_out;
  wire [63:0] cout_drain_IO_L1_out_wrapper408_U0_fifo_cout_drain_out_V_V_din_pass_1_in;
  wire fifo_cout_drain_cout_drain_IO_L1_out_2_6_V_V_full_n_pass_1_out;
  wire cout_drain_IO_L1_out_wrapper408_U0_fifo_cout_drain_out_V_V_write_pass_1_in;
  wire [255:0] PE_wrapper213_U0_fifo_w_out_V_V_din_pass_0_out;
  wire fifo_w_PE_5_4_V_V_full_n_pass_0_in;
  wire PE_wrapper213_U0_fifo_w_out_V_V_write_pass_0_out;
  wire [63:0] cout_drain_IO_L2_out568_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  wire fifo_cout_drain_cout_drain_IO_L2_out_0_V_V_full_n_pass_0_in;
  wire cout_drain_IO_L2_out568_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  wire [31:0] PE_wrapper176_U0_fifo_cout_drain_out_V_din_pass_1_in;
  wire fifo_cout_drain_PE_2_2_V_full_n_pass_1_out;
  wire PE_wrapper176_U0_fifo_cout_drain_out_V_write_pass_1_in;
  wire ap_start_Boundary_X6Y0_To_X6Y2_in;
  wire ap_rst_n_Boundary_X6Y0_To_X6Y2_in;
  wire ap_done_Boundary_X6Y0_To_X6Y2_out;
  wire ap_start_Boundary_X6Y2_To_X8Y2_out;
  wire ap_rst_n_Boundary_X6Y2_To_X8Y2_out;
  wire ap_done_Boundary_X6Y2_To_X8Y2_in;
  wire [63:0] cout_drain_IO_L2_out564_U0_fifo_cout_drain_out_V_V_din_pass_0_in;
  wire [63:0] cout_drain_IO_L2_out564_U0_fifo_cout_drain_out_V_V_din_pass_1_out;
  wire fifo_cout_drain_cout_drain_IO_L2_out_4_V_V_full_n_pass_0_out;
  wire fifo_cout_drain_cout_drain_IO_L2_out_4_V_V_full_n_pass_1_in;
  wire cout_drain_IO_L2_out564_U0_fifo_cout_drain_out_V_V_write_pass_0_in;
  wire cout_drain_IO_L2_out564_U0_fifo_cout_drain_out_V_V_write_pass_1_out;
  wire [31:0] PE_wrapper165_U0_fifo_cout_drain_out_V_din_pass_0_in;
  wire [31:0] PE_wrapper165_U0_fifo_cout_drain_out_V_din_pass_1_out;
  wire fifo_cout_drain_PE_1_3_V_full_n_pass_0_out;
  wire fifo_cout_drain_PE_1_3_V_full_n_pass_1_in;
  wire PE_wrapper165_U0_fifo_cout_drain_out_V_write_pass_0_in;
  wire PE_wrapper165_U0_fifo_cout_drain_out_V_write_pass_1_out;
  wire [31:0] PE_wrapper153_U0_fifo_cout_drain_out_V_din_pass_0_in;
  wire [31:0] PE_wrapper153_U0_fifo_cout_drain_out_V_din_pass_1_out;
  wire fifo_cout_drain_PE_0_3_V_full_n_pass_0_out;
  wire fifo_cout_drain_PE_0_3_V_full_n_pass_1_in;
  wire PE_wrapper153_U0_fifo_cout_drain_out_V_write_pass_0_in;
  wire PE_wrapper153_U0_fifo_cout_drain_out_V_write_pass_1_out;
  wire [31:0] PE_wrapper177_U0_fifo_cout_drain_out_V_din_pass_0_in;
  wire [31:0] PE_wrapper177_U0_fifo_cout_drain_out_V_din_pass_1_out;
  wire fifo_cout_drain_PE_2_3_V_full_n_pass_0_out;
  wire fifo_cout_drain_PE_2_3_V_full_n_pass_1_in;
  wire PE_wrapper177_U0_fifo_cout_drain_out_V_write_pass_0_in;
  wire PE_wrapper177_U0_fifo_cout_drain_out_V_write_pass_1_out;
  wire [31:0] PE_wrapper164_U0_fifo_cout_drain_out_V_din_pass_0_in;
  wire [31:0] PE_wrapper164_U0_fifo_cout_drain_out_V_din_pass_1_out;
  wire fifo_cout_drain_PE_1_2_V_full_n_pass_0_out;
  wire fifo_cout_drain_PE_1_2_V_full_n_pass_1_in;
  wire PE_wrapper164_U0_fifo_cout_drain_out_V_write_pass_0_in;
  wire PE_wrapper164_U0_fifo_cout_drain_out_V_write_pass_1_out;
  wire [31:0] PE_wrapper189_U0_fifo_cout_drain_out_V_din_pass_0_in;
  wire [31:0] PE_wrapper189_U0_fifo_cout_drain_out_V_din_pass_1_out;
  wire fifo_cout_drain_PE_3_3_V_full_n_pass_0_out;
  wire fifo_cout_drain_PE_3_3_V_full_n_pass_1_in;
  wire PE_wrapper189_U0_fifo_cout_drain_out_V_write_pass_0_in;
  wire PE_wrapper189_U0_fifo_cout_drain_out_V_write_pass_1_out;
  wire [31:0] PE_wrapper152_U0_fifo_cout_drain_out_V_din_pass_0_in;
  wire [31:0] PE_wrapper152_U0_fifo_cout_drain_out_V_din_pass_1_out;
  wire fifo_cout_drain_PE_0_2_V_full_n_pass_0_out;
  wire fifo_cout_drain_PE_0_2_V_full_n_pass_1_in;
  wire PE_wrapper152_U0_fifo_cout_drain_out_V_write_pass_0_in;
  wire PE_wrapper152_U0_fifo_cout_drain_out_V_write_pass_1_out;
  wire [31:0] PE_wrapper176_U0_fifo_cout_drain_out_V_din_pass_0_in;
  wire [31:0] PE_wrapper176_U0_fifo_cout_drain_out_V_din_pass_1_out;
  wire fifo_cout_drain_PE_2_2_V_full_n_pass_0_out;
  wire fifo_cout_drain_PE_2_2_V_full_n_pass_1_in;
  wire PE_wrapper176_U0_fifo_cout_drain_out_V_write_pass_0_in;
  wire PE_wrapper176_U0_fifo_cout_drain_out_V_write_pass_1_out;
  wire [255:0] PE_wrapper165_U0_fifo_w_out_V_V_din_pass_0_in;
  wire [255:0] PE_wrapper165_U0_fifo_w_out_V_V_din_pass_1_out;
  wire fifo_w_PE_1_4_V_V_full_n_pass_0_out;
  wire fifo_w_PE_1_4_V_V_full_n_pass_1_in;
  wire PE_wrapper165_U0_fifo_w_out_V_V_write_pass_0_in;
  wire PE_wrapper165_U0_fifo_w_out_V_V_write_pass_1_out;
  wire [255:0] cin_IO_L2_in127_U0_fifo_cin_out_V_V_din_pass_0_in;
  wire [255:0] cin_IO_L2_in127_U0_fifo_cin_out_V_V_din_pass_1_out;
  wire fifo_cin_cin_IO_L2_in_4_V_V_full_n_pass_0_out;
  wire fifo_cin_cin_IO_L2_in_4_V_V_full_n_pass_1_in;
  wire cin_IO_L2_in127_U0_fifo_cin_out_V_V_write_pass_0_in;
  wire cin_IO_L2_in127_U0_fifo_cin_out_V_V_write_pass_1_out;
  wire [255:0] PE_wrapper177_U0_fifo_w_out_V_V_din_pass_0_in;
  wire [255:0] PE_wrapper177_U0_fifo_w_out_V_V_din_pass_1_out;
  wire fifo_w_PE_2_4_V_V_full_n_pass_0_out;
  wire fifo_w_PE_2_4_V_V_full_n_pass_1_in;
  wire PE_wrapper177_U0_fifo_w_out_V_V_write_pass_0_in;
  wire PE_wrapper177_U0_fifo_w_out_V_V_write_pass_1_out;
  wire [255:0] PE_wrapper153_U0_fifo_w_out_V_V_din_pass_0_in;
  wire [255:0] PE_wrapper153_U0_fifo_w_out_V_V_din_pass_1_out;
  wire fifo_w_PE_0_4_V_V_full_n_pass_0_out;
  wire fifo_w_PE_0_4_V_V_full_n_pass_1_in;
  wire PE_wrapper153_U0_fifo_w_out_V_V_write_pass_0_in;
  wire PE_wrapper153_U0_fifo_w_out_V_V_write_pass_1_out;
  wire [255:0] PE_wrapper189_U0_fifo_w_out_V_V_din_pass_0_in;
  wire [255:0] PE_wrapper189_U0_fifo_w_out_V_V_din_pass_1_out;
  wire fifo_w_PE_3_4_V_V_full_n_pass_0_out;
  wire fifo_w_PE_3_4_V_V_full_n_pass_1_in;
  wire PE_wrapper189_U0_fifo_w_out_V_V_write_pass_0_in;
  wire PE_wrapper189_U0_fifo_w_out_V_V_write_pass_1_out;
  wire [63:0] cout_drain_IO_L2_out568_U0_fifo_cout_drain_out_V_V_din_pass_0_in;
  wire [63:0] cout_drain_IO_L2_out568_U0_fifo_cout_drain_out_V_V_din_pass_1_out;
  wire fifo_cout_drain_cout_drain_IO_L2_out_0_V_V_full_n_pass_0_out;
  wire fifo_cout_drain_cout_drain_IO_L2_out_0_V_V_full_n_pass_1_in;
  wire cout_drain_IO_L2_out568_U0_fifo_cout_drain_out_V_V_write_pass_0_in;
  wire cout_drain_IO_L2_out568_U0_fifo_cout_drain_out_V_V_write_pass_1_out;
  wire [255:0] w_IO_L2_in140_U0_fifo_w_out_V_V_din_pass_0_out;
  wire fifo_w_w_IO_L2_in_6_V_V_full_n_pass_0_in;
  wire w_IO_L2_in140_U0_fifo_w_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper187_U0_fifo_w_out_V_V_din_pass_1_in;
  wire fifo_w_PE_3_2_V_V_full_n_pass_1_out;
  wire PE_wrapper187_U0_fifo_w_out_V_V_write_pass_1_in;
  wire [255:0] PE_wrapper188_U0_fifo_w_out_V_V_din_pass_0_out;
  wire fifo_w_PE_3_3_V_V_full_n_pass_0_in;
  wire PE_wrapper188_U0_fifo_w_out_V_V_write_pass_0_out;
  wire [31:0] PE_wrapper200_U0_fifo_cout_drain_out_V_din_pass_0_out;
  wire fifo_cout_drain_PE_4_2_V_full_n_pass_0_in;
  wire PE_wrapper200_U0_fifo_cout_drain_out_V_write_pass_0_out;
  wire [31:0] PE_wrapper188_U0_fifo_cout_drain_out_V_din_pass_0_out;
  wire fifo_cout_drain_PE_3_2_V_full_n_pass_0_in;
  wire PE_wrapper188_U0_fifo_cout_drain_out_V_write_pass_0_out;
  wire [255:0] PE_wrapper210_U0_fifo_w_out_V_V_din_pass_0_out;
  wire fifo_w_PE_5_1_V_V_full_n_pass_0_in;
  wire PE_wrapper210_U0_fifo_w_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper201_U0_fifo_cin_out_V_V_din_pass_0_out;
  wire fifo_cin_PE_5_3_V_V_full_n_pass_0_in;
  wire PE_wrapper201_U0_fifo_cin_out_V_V_write_pass_0_out;
  wire [63:0] cout_drain_IO_L1_out_wrapper398_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_1_0_V_V_full_n_pass_0_in;
  wire cout_drain_IO_L1_out_wrapper398_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper199_U0_fifo_cin_out_V_V_din_pass_0_out;
  wire fifo_cin_PE_5_1_V_V_full_n_pass_0_in;
  wire PE_wrapper199_U0_fifo_cin_out_V_V_write_pass_0_out;
  wire [31:0] PE_wrapper163_U0_fifo_cout_drain_out_V_din_pass_1_in;
  wire fifo_cout_drain_PE_1_1_V_full_n_pass_1_out;
  wire PE_wrapper163_U0_fifo_cout_drain_out_V_write_pass_1_in;
  wire [31:0] PE_wrapper211_U0_fifo_cout_drain_out_V_din_pass_0_in;
  wire fifo_cout_drain_PE_5_1_V_full_n_pass_0_out;
  wire PE_wrapper211_U0_fifo_cout_drain_out_V_write_pass_0_in;
  wire [63:0] cout_drain_IO_L1_out_wrapper378_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_0_4_V_V_full_n_pass_0_in;
  wire cout_drain_IO_L1_out_wrapper378_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  wire [31:0] PE_wrapper175_U0_fifo_cout_drain_out_V_din_pass_1_in;
  wire fifo_cout_drain_PE_2_1_V_full_n_pass_1_out;
  wire PE_wrapper175_U0_fifo_cout_drain_out_V_write_pass_1_in;
  wire [31:0] PE_wrapper201_U0_fifo_cout_drain_out_V_din_pass_0_out;
  wire fifo_cout_drain_PE_4_3_V_full_n_pass_0_in;
  wire PE_wrapper201_U0_fifo_cout_drain_out_V_write_pass_0_out;
  wire [255:0] PE_wrapper187_U0_fifo_cin_out_V_V_din_pass_1_in;
  wire fifo_cin_PE_4_1_V_V_full_n_pass_1_out;
  wire PE_wrapper187_U0_fifo_cin_out_V_V_write_pass_1_in;
  wire [255:0] PE_wrapper186_U0_fifo_cin_out_V_V_din_pass_1_in;
  wire fifo_cin_PE_4_0_V_V_full_n_pass_1_out;
  wire PE_wrapper186_U0_fifo_cin_out_V_V_write_pass_1_in;
  wire [255:0] PE_wrapper201_U0_fifo_w_out_V_V_din_pass_0_out;
  wire fifo_w_PE_4_4_V_V_full_n_pass_0_in;
  wire PE_wrapper201_U0_fifo_w_out_V_V_write_pass_0_out;
  wire [31:0] PE_wrapper187_U0_fifo_cout_drain_out_V_din_pass_1_in;
  wire fifo_cout_drain_PE_3_1_V_full_n_pass_1_out;
  wire PE_wrapper187_U0_fifo_cout_drain_out_V_write_pass_1_in;
  wire [255:0] w_IO_L2_in137_U0_fifo_w_out_V_V_din_pass_1_in;
  wire fifo_w_w_IO_L2_in_3_V_V_full_n_pass_1_out;
  wire w_IO_L2_in137_U0_fifo_w_out_V_V_write_pass_1_in;
  wire [63:0] cout_drain_IO_L1_out_wrapper376_U0_fifo_cout_drain_out_V_V_din_pass_2_in;
  wire fifo_cout_drain_cout_drain_IO_L1_out_0_6_V_V_full_n_pass_2_out;
  wire cout_drain_IO_L1_out_wrapper376_U0_fifo_cout_drain_out_V_V_write_pass_2_in;
  wire [31:0] PE_wrapper151_U0_fifo_cout_drain_out_V_din_pass_1_in;
  wire fifo_cout_drain_PE_0_1_V_full_n_pass_1_out;
  wire PE_wrapper151_U0_fifo_cout_drain_out_V_write_pass_1_in;
  wire [255:0] w_IO_L2_in138_U0_fifo_w_local_out_V_V_din_pass_0_out;
  wire fifo_w_PE_3_0_V_V_full_n_pass_0_in;
  wire w_IO_L2_in138_U0_fifo_w_local_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper200_U0_fifo_cin_out_V_V_din_pass_0_out;
  wire fifo_cin_PE_5_2_V_V_full_n_pass_0_in;
  wire PE_wrapper200_U0_fifo_cin_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper189_U0_fifo_cin_out_V_V_din_pass_0_in;
  wire fifo_cin_PE_4_3_V_V_full_n_pass_0_out;
  wire PE_wrapper189_U0_fifo_cin_out_V_V_write_pass_0_in;
  wire [255:0] PE_wrapper176_U0_fifo_cin_out_V_V_din_pass_0_in;
  wire fifo_cin_PE_3_2_V_V_full_n_pass_0_out;
  wire PE_wrapper176_U0_fifo_cin_out_V_V_write_pass_0_in;
  wire [255:0] PE_wrapper210_U0_fifo_cin_out_V_V_din_pass_0_out;
  wire fifo_cin_PE_6_0_V_V_full_n_pass_0_in;
  wire PE_wrapper210_U0_fifo_cin_out_V_V_write_pass_0_out;
  wire [63:0] cout_drain_IO_L1_out_wrapper392_U0_fifo_cout_drain_out_V_V_din_pass_2_in;
  wire fifo_cout_drain_cout_drain_IO_L1_out_1_6_V_V_full_n_pass_2_out;
  wire cout_drain_IO_L1_out_wrapper392_U0_fifo_cout_drain_out_V_V_write_pass_2_in;
  wire ap_start_Boundary_X6Y2_To_X8Y2_in;
  wire ap_rst_n_Boundary_X6Y2_To_X8Y2_in;
  wire ap_done_Boundary_X6Y2_To_X8Y2_out;
  wire ap_start_Boundary_X6Y4_To_X8Y4_out;
  wire ap_rst_n_Boundary_X6Y4_To_X8Y4_out;
  wire ap_done_Boundary_X6Y4_To_X8Y4_in;
  wire [255:0] PE_wrapper214_U0_fifo_w_out_V_V_din_pass_0_in;
  wire [255:0] PE_wrapper214_U0_fifo_w_out_V_V_din_pass_1_out;
  wire fifo_w_PE_5_5_V_V_full_n_pass_0_out;
  wire fifo_w_PE_5_5_V_V_full_n_pass_1_in;
  wire PE_wrapper214_U0_fifo_w_out_V_V_write_pass_0_in;
  wire PE_wrapper214_U0_fifo_w_out_V_V_write_pass_1_out;
  wire [255:0] PE_wrapper202_U0_fifo_w_out_V_V_din_pass_0_in;
  wire [255:0] PE_wrapper202_U0_fifo_w_out_V_V_din_pass_1_out;
  wire fifo_w_PE_4_5_V_V_full_n_pass_0_out;
  wire fifo_w_PE_4_5_V_V_full_n_pass_1_in;
  wire PE_wrapper202_U0_fifo_w_out_V_V_write_pass_0_in;
  wire PE_wrapper202_U0_fifo_w_out_V_V_write_pass_1_out;
  wire [63:0] kernel0_entry12_U0_cout_V_out_din_pass_2_in;
  wire [63:0] kernel0_entry12_U0_cout_V_out_din_pass_3_out;
  wire cout_V_c_full_n_pass_2_out;
  wire cout_V_c_full_n_pass_3_in;
  wire kernel0_entry12_U0_cout_V_out_write_pass_2_in;
  wire kernel0_entry12_U0_cout_V_out_write_pass_3_out;
  wire [255:0] PE_wrapper243_U0_fifo_w_out_V_V_din_pass_0_in;
  wire [255:0] PE_wrapper243_U0_fifo_w_out_V_V_din_pass_1_out;
  wire fifo_w_PE_7_10_V_V_full_n_pass_0_out;
  wire fifo_w_PE_7_10_V_V_full_n_pass_1_in;
  wire PE_wrapper243_U0_fifo_w_out_V_V_write_pass_0_in;
  wire PE_wrapper243_U0_fifo_w_out_V_V_write_pass_1_out;
  wire [31:0] PE_wrapper243_U0_fifo_cout_drain_out_V_din_pass_0_in;
  wire [31:0] PE_wrapper243_U0_fifo_cout_drain_out_V_din_pass_1_out;
  wire fifo_cout_drain_PE_7_9_V_full_n_pass_0_out;
  wire fifo_cout_drain_PE_7_9_V_full_n_pass_1_in;
  wire PE_wrapper243_U0_fifo_cout_drain_out_V_write_pass_0_in;
  wire PE_wrapper243_U0_fifo_cout_drain_out_V_write_pass_1_out;
  wire [255:0] PE_wrapper243_U0_fifo_cin_out_V_V_din_pass_0_in;
  wire [255:0] PE_wrapper243_U0_fifo_cin_out_V_V_din_pass_1_out;
  wire fifo_cin_PE_8_9_V_V_full_n_pass_0_out;
  wire fifo_cin_PE_8_9_V_V_full_n_pass_1_in;
  wire PE_wrapper243_U0_fifo_cin_out_V_V_write_pass_0_in;
  wire PE_wrapper243_U0_fifo_cin_out_V_V_write_pass_1_out;
  wire [255:0] PE_wrapper191_U0_fifo_cin_out_V_V_din_pass_0_out;
  wire fifo_cin_PE_4_5_V_V_full_n_pass_0_in;
  wire PE_wrapper191_U0_fifo_cin_out_V_V_write_pass_0_out;
  wire [31:0] PE_wrapper191_U0_fifo_cout_drain_out_V_din_pass_0_out;
  wire fifo_cout_drain_PE_3_5_V_full_n_pass_0_in;
  wire PE_wrapper191_U0_fifo_cout_drain_out_V_write_pass_0_out;
  wire [255:0] PE_wrapper192_U0_fifo_cin_out_V_V_din_pass_0_out;
  wire fifo_cin_PE_4_6_V_V_full_n_pass_0_in;
  wire PE_wrapper192_U0_fifo_cin_out_V_V_write_pass_0_out;
  wire [31:0] PE_wrapper192_U0_fifo_cout_drain_out_V_din_pass_0_out;
  wire fifo_cout_drain_PE_3_6_V_full_n_pass_0_in;
  wire PE_wrapper192_U0_fifo_cout_drain_out_V_write_pass_0_out;
  wire [255:0] PE_wrapper192_U0_fifo_w_out_V_V_din_pass_0_out;
  wire fifo_w_PE_3_7_V_V_full_n_pass_0_in;
  wire PE_wrapper192_U0_fifo_w_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper190_U0_fifo_w_out_V_V_din_pass_1_in;
  wire fifo_w_PE_3_5_V_V_full_n_pass_1_out;
  wire PE_wrapper190_U0_fifo_w_out_V_V_write_pass_1_in;
  wire [255:0] PE_wrapper179_U0_fifo_cin_out_V_V_din_pass_1_in;
  wire fifo_cin_PE_3_5_V_V_full_n_pass_1_out;
  wire PE_wrapper179_U0_fifo_cin_out_V_V_write_pass_1_in;
  wire [255:0] PE_wrapper180_U0_fifo_cin_out_V_V_din_pass_0_in;
  wire fifo_cin_PE_3_6_V_V_full_n_pass_0_out;
  wire PE_wrapper180_U0_fifo_cin_out_V_V_write_pass_0_in;
  wire ap_start_Boundary_X4Y6_To_X6Y6_in;
  wire ap_rst_n_Boundary_X4Y6_To_X6Y6_in;
  wire ap_done_Boundary_X4Y6_To_X6Y6_out;
  wire ap_start_Boundary_X4Y8_To_X6Y8_out;
  wire ap_rst_n_Boundary_X4Y8_To_X6Y8_out;
  wire ap_done_Boundary_X4Y8_To_X6Y8_in;
  wire [63:0] cout_drain_IO_L2_out568_U0_fifo_cout_drain_out_V_V_din_pass_1_in;
  wire [63:0] cout_drain_IO_L2_out568_U0_fifo_cout_drain_out_V_V_din_pass_2_out;
  wire fifo_cout_drain_cout_drain_IO_L2_out_0_V_V_full_n_pass_1_out;
  wire fifo_cout_drain_cout_drain_IO_L2_out_0_V_V_full_n_pass_2_in;
  wire cout_drain_IO_L2_out568_U0_fifo_cout_drain_out_V_V_write_pass_1_in;
  wire cout_drain_IO_L2_out568_U0_fifo_cout_drain_out_V_V_write_pass_2_out;
  wire [255:0] PE_wrapper165_U0_fifo_w_out_V_V_din_pass_1_in;
  wire fifo_w_PE_1_4_V_V_full_n_pass_1_out;
  wire PE_wrapper165_U0_fifo_w_out_V_V_write_pass_1_in;
  wire [63:0] cout_drain_IO_L2_out564_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  wire fifo_cout_drain_cout_drain_IO_L2_out_4_V_V_full_n_pass_0_in;
  wire cout_drain_IO_L2_out564_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  wire [255:0] cin_IO_L2_in127_U0_fifo_cin_out_V_V_din_pass_1_in;
  wire fifo_cin_cin_IO_L2_in_4_V_V_full_n_pass_1_out;
  wire cin_IO_L2_in127_U0_fifo_cin_out_V_V_write_pass_1_in;
  wire [255:0] PE_wrapper179_U0_fifo_w_out_V_V_din_pass_0_out;
  wire fifo_w_PE_2_6_V_V_full_n_pass_0_in;
  wire PE_wrapper179_U0_fifo_w_out_V_V_write_pass_0_out;
  wire [255:0] cin_IO_L2_in128_U0_fifo_cin_out_V_V_din_pass_0_out;
  wire fifo_cin_cin_IO_L2_in_5_V_V_full_n_pass_0_in;
  wire cin_IO_L2_in128_U0_fifo_cin_out_V_V_write_pass_0_out;
  wire [31:0] PE_wrapper179_U0_fifo_cout_drain_out_V_din_pass_0_out;
  wire fifo_cout_drain_PE_2_5_V_full_n_pass_0_in;
  wire PE_wrapper179_U0_fifo_cout_drain_out_V_write_pass_0_out;
  wire [255:0] PE_wrapper177_U0_fifo_w_out_V_V_din_pass_1_in;
  wire fifo_w_PE_2_4_V_V_full_n_pass_1_out;
  wire PE_wrapper177_U0_fifo_w_out_V_V_write_pass_1_in;
  wire [255:0] PE_wrapper153_U0_fifo_w_out_V_V_din_pass_1_in;
  wire fifo_w_PE_0_4_V_V_full_n_pass_1_out;
  wire PE_wrapper153_U0_fifo_w_out_V_V_write_pass_1_in;
  wire [255:0] PE_wrapper190_U0_fifo_cin_out_V_V_din_pass_0_out;
  wire fifo_cin_PE_4_4_V_V_full_n_pass_0_in;
  wire PE_wrapper190_U0_fifo_cin_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper166_U0_fifo_w_out_V_V_din_pass_0_out;
  wire fifo_w_PE_1_5_V_V_full_n_pass_0_in;
  wire PE_wrapper166_U0_fifo_w_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper154_U0_fifo_w_out_V_V_din_pass_0_out;
  wire fifo_w_PE_0_5_V_V_full_n_pass_0_in;
  wire PE_wrapper154_U0_fifo_w_out_V_V_write_pass_0_out;
  wire [63:0] cout_drain_IO_L2_out563_U0_fifo_cout_drain_out_V_V_din_pass_0_in;
  wire fifo_cout_drain_cout_drain_IO_L2_out_5_V_V_full_n_pass_0_out;
  wire cout_drain_IO_L2_out563_U0_fifo_cout_drain_out_V_V_write_pass_0_in;
  wire [255:0] PE_wrapper190_U0_fifo_w_out_V_V_din_pass_0_out;
  wire fifo_w_PE_3_5_V_V_full_n_pass_0_in;
  wire PE_wrapper190_U0_fifo_w_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper179_U0_fifo_cin_out_V_V_din_pass_0_out;
  wire fifo_cin_PE_3_5_V_V_full_n_pass_0_in;
  wire PE_wrapper179_U0_fifo_cin_out_V_V_write_pass_0_out;
  wire [31:0] PE_wrapper202_U0_fifo_cout_drain_out_V_din_pass_0_in;
  wire fifo_cout_drain_PE_4_4_V_full_n_pass_0_out;
  wire PE_wrapper202_U0_fifo_cout_drain_out_V_write_pass_0_in;
  wire [255:0] PE_wrapper189_U0_fifo_w_out_V_V_din_pass_1_in;
  wire fifo_w_PE_3_4_V_V_full_n_pass_1_out;
  wire PE_wrapper189_U0_fifo_w_out_V_V_write_pass_1_in;
  wire [255:0] PE_wrapper167_U0_fifo_cin_out_V_V_din_pass_0_in;
  wire fifo_cin_PE_2_5_V_V_full_n_pass_0_out;
  wire PE_wrapper167_U0_fifo_cin_out_V_V_write_pass_0_in;
  wire [63:0] cout_drain_IO_L1_out_wrapper441_U0_fifo_cout_drain_out_V_V_din_pass_0_in;
  wire fifo_cout_drain_cout_drain_IO_L1_out_4_5_V_V_full_n_pass_0_out;
  wire cout_drain_IO_L1_out_wrapper441_U0_fifo_cout_drain_out_V_V_write_pass_0_in;
  wire ap_start_Boundary_X6Y4_To_X8Y4_in;
  wire ap_rst_n_Boundary_X6Y4_To_X8Y4_in;
  wire ap_done_Boundary_X6Y4_To_X8Y4_out;
  wire ap_start_Boundary_X6Y6_To_X8Y6_out;
  wire ap_rst_n_Boundary_X6Y6_To_X8Y6_out;
  wire ap_done_Boundary_X6Y6_To_X8Y6_in;
  wire [255:0] PE_wrapper192_U0_fifo_w_out_V_V_din_pass_0_in;
  wire [255:0] PE_wrapper192_U0_fifo_w_out_V_V_din_pass_1_out;
  wire fifo_w_PE_3_7_V_V_full_n_pass_0_out;
  wire fifo_w_PE_3_7_V_V_full_n_pass_1_in;
  wire PE_wrapper192_U0_fifo_w_out_V_V_write_pass_0_in;
  wire PE_wrapper192_U0_fifo_w_out_V_V_write_pass_1_out;
  wire [63:0] cout_drain_IO_L2_out568_U0_fifo_cout_drain_out_V_V_din_pass_2_in;
  wire [63:0] cout_drain_IO_L2_out568_U0_fifo_cout_drain_out_V_V_din_pass_3_out;
  wire fifo_cout_drain_cout_drain_IO_L2_out_0_V_V_full_n_pass_2_out;
  wire fifo_cout_drain_cout_drain_IO_L2_out_0_V_V_full_n_pass_3_in;
  wire cout_drain_IO_L2_out568_U0_fifo_cout_drain_out_V_V_write_pass_2_in;
  wire cout_drain_IO_L2_out568_U0_fifo_cout_drain_out_V_V_write_pass_3_out;
  wire [255:0] PE_wrapper168_U0_fifo_w_out_V_V_din_pass_0_out;
  wire fifo_w_PE_1_7_V_V_full_n_pass_0_in;
  wire PE_wrapper168_U0_fifo_w_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper179_U0_fifo_w_out_V_V_din_pass_0_in;
  wire fifo_w_PE_2_6_V_V_full_n_pass_0_out;
  wire PE_wrapper179_U0_fifo_w_out_V_V_write_pass_0_in;
  wire [255:0] cin_IO_L2_in128_U0_fifo_cin_out_V_V_din_pass_0_in;
  wire fifo_cin_cin_IO_L2_in_5_V_V_full_n_pass_0_out;
  wire cin_IO_L2_in128_U0_fifo_cin_out_V_V_write_pass_0_in;
  wire [63:0] cout_drain_IO_L2_out561_U0_fifo_cout_drain_out_V_V_din_pass_0_in;
  wire fifo_cout_drain_cout_drain_IO_L2_out_7_V_V_full_n_pass_0_out;
  wire cout_drain_IO_L2_out561_U0_fifo_cout_drain_out_V_V_write_pass_0_in;
  wire [255:0] PE_wrapper242_U0_fifo_w_out_V_V_din_pass_2_in;
  wire fifo_w_PE_7_9_V_V_full_n_pass_2_out;
  wire PE_wrapper242_U0_fifo_w_out_V_V_write_pass_2_in;
  wire [31:0] PE_wrapper179_U0_fifo_cout_drain_out_V_din_pass_0_in;
  wire fifo_cout_drain_PE_2_5_V_full_n_pass_0_out;
  wire PE_wrapper179_U0_fifo_cout_drain_out_V_write_pass_0_in;
  wire [255:0] cin_IO_L2_in130_U0_fifo_cin_out_V_V_din_pass_0_out;
  wire fifo_cin_cin_IO_L2_in_7_V_V_full_n_pass_0_in;
  wire cin_IO_L2_in130_U0_fifo_cin_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper166_U0_fifo_w_out_V_V_din_pass_0_in;
  wire fifo_w_PE_1_5_V_V_full_n_pass_0_out;
  wire PE_wrapper166_U0_fifo_w_out_V_V_write_pass_0_in;
  wire [255:0] PE_wrapper243_U0_fifo_w_out_V_V_din_pass_0_out;
  wire fifo_w_PE_7_10_V_V_full_n_pass_0_in;
  wire PE_wrapper243_U0_fifo_w_out_V_V_write_pass_0_out;
  wire [31:0] PE_wrapper243_U0_fifo_cout_drain_out_V_din_pass_0_out;
  wire fifo_cout_drain_PE_7_9_V_full_n_pass_0_in;
  wire PE_wrapper243_U0_fifo_cout_drain_out_V_write_pass_0_out;
  wire [255:0] PE_wrapper243_U0_fifo_cin_out_V_V_din_pass_0_out;
  wire fifo_cin_PE_8_9_V_V_full_n_pass_0_in;
  wire PE_wrapper243_U0_fifo_cin_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper154_U0_fifo_w_out_V_V_din_pass_0_in;
  wire fifo_w_PE_0_5_V_V_full_n_pass_0_out;
  wire PE_wrapper154_U0_fifo_w_out_V_V_write_pass_0_in;
  wire [255:0] PE_wrapper156_U0_fifo_w_out_V_V_din_pass_0_out;
  wire fifo_w_PE_0_7_V_V_full_n_pass_0_in;
  wire PE_wrapper156_U0_fifo_w_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper180_U0_fifo_cin_out_V_V_din_pass_0_out;
  wire fifo_cin_PE_3_6_V_V_full_n_pass_0_in;
  wire PE_wrapper180_U0_fifo_cin_out_V_V_write_pass_0_out;
  wire [63:0] cout_drain_IO_L2_out563_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  wire fifo_cout_drain_cout_drain_IO_L2_out_5_V_V_full_n_pass_0_in;
  wire cout_drain_IO_L2_out563_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  wire [31:0] PE_wrapper191_U0_fifo_cout_drain_out_V_din_pass_0_in;
  wire fifo_cout_drain_PE_3_5_V_full_n_pass_0_out;
  wire PE_wrapper191_U0_fifo_cout_drain_out_V_write_pass_0_in;
  wire [63:0] cout_drain_IO_L1_out_wrapper474_U0_fifo_cout_drain_out_V_V_din_pass_1_in;
  wire fifo_cout_drain_cout_drain_IO_L1_out_6_4_V_V_full_n_pass_1_out;
  wire cout_drain_IO_L1_out_wrapper474_U0_fifo_cout_drain_out_V_V_write_pass_1_in;
  wire [63:0] cout_drain_IO_L1_out_wrapper458_U0_fifo_cout_drain_out_V_V_din_pass_1_in;
  wire fifo_cout_drain_cout_drain_IO_L1_out_5_4_V_V_full_n_pass_1_out;
  wire cout_drain_IO_L1_out_wrapper458_U0_fifo_cout_drain_out_V_V_write_pass_1_in;
  wire [255:0] PE_wrapper180_U0_fifo_w_out_V_V_din_pass_0_out;
  wire fifo_w_PE_2_7_V_V_full_n_pass_0_in;
  wire PE_wrapper180_U0_fifo_w_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper167_U0_fifo_cin_out_V_V_din_pass_0_out;
  wire fifo_cin_PE_2_5_V_V_full_n_pass_0_in;
  wire PE_wrapper167_U0_fifo_cin_out_V_V_write_pass_0_out;
  wire [31:0] PE_wrapper192_U0_fifo_cout_drain_out_V_din_pass_0_in;
  wire fifo_cout_drain_PE_3_6_V_full_n_pass_0_out;
  wire PE_wrapper192_U0_fifo_cout_drain_out_V_write_pass_0_in;
  wire [255:0] PE_wrapper231_U0_fifo_cin_out_V_V_din_pass_4_in;
  wire fifo_cin_PE_7_9_V_V_full_n_pass_4_out;
  wire PE_wrapper231_U0_fifo_cin_out_V_V_write_pass_4_in;
  wire ap_start_Boundary_X6Y6_To_X8Y6_in;
  wire ap_rst_n_Boundary_X6Y6_To_X8Y6_in;
  wire ap_done_Boundary_X6Y6_To_X8Y6_out;
  wire ap_start_Boundary_X6Y8_To_X8Y8_out;
  wire ap_rst_n_Boundary_X6Y8_To_X8Y8_out;
  wire ap_done_Boundary_X6Y8_To_X8Y8_in;
  wire [255:0] PE_wrapper251_U0_fifo_w_out_V_V_din_pass_0_in;
  wire [255:0] PE_wrapper251_U0_fifo_w_out_V_V_din_pass_1_out;
  wire fifo_w_PE_8_6_V_V_full_n_pass_0_out;
  wire fifo_w_PE_8_6_V_V_full_n_pass_1_in;
  wire PE_wrapper251_U0_fifo_w_out_V_V_write_pass_0_in;
  wire PE_wrapper251_U0_fifo_w_out_V_V_write_pass_1_out;
  wire [255:0] PE_wrapper239_U0_fifo_w_out_V_V_din_pass_0_in;
  wire [255:0] PE_wrapper239_U0_fifo_w_out_V_V_din_pass_1_out;
  wire fifo_w_PE_7_6_V_V_full_n_pass_0_out;
  wire fifo_w_PE_7_6_V_V_full_n_pass_1_in;
  wire PE_wrapper239_U0_fifo_w_out_V_V_write_pass_0_in;
  wire PE_wrapper239_U0_fifo_w_out_V_V_write_pass_1_out;
  wire [63:0] cout_drain_IO_L1_out_wrapper469_U0_fifo_cout_drain_out_V_V_din_pass_0_in;
  wire [63:0] cout_drain_IO_L1_out_wrapper469_U0_fifo_cout_drain_out_V_V_din_pass_1_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_6_9_V_V_full_n_pass_0_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_6_9_V_V_full_n_pass_1_in;
  wire cout_drain_IO_L1_out_wrapper469_U0_fifo_cout_drain_out_V_V_write_pass_0_in;
  wire cout_drain_IO_L1_out_wrapper469_U0_fifo_cout_drain_out_V_V_write_pass_1_out;
  wire [63:0] kernel0_entry12_U0_cout_V_out_din_pass_3_in;
  wire [63:0] kernel0_entry12_U0_cout_V_out_din_pass_4_out;
  wire cout_V_c_full_n_pass_3_out;
  wire cout_V_c_full_n_pass_4_in;
  wire kernel0_entry12_U0_cout_V_out_write_pass_3_in;
  wire kernel0_entry12_U0_cout_V_out_write_pass_4_out;
  wire [255:0] PE_wrapper243_U0_fifo_w_out_V_V_din_pass_1_in;
  wire [255:0] PE_wrapper243_U0_fifo_w_out_V_V_din_pass_2_out;
  wire fifo_w_PE_7_10_V_V_full_n_pass_1_out;
  wire fifo_w_PE_7_10_V_V_full_n_pass_2_in;
  wire PE_wrapper243_U0_fifo_w_out_V_V_write_pass_1_in;
  wire PE_wrapper243_U0_fifo_w_out_V_V_write_pass_2_out;
  wire [31:0] PE_wrapper243_U0_fifo_cout_drain_out_V_din_pass_1_in;
  wire [31:0] PE_wrapper243_U0_fifo_cout_drain_out_V_din_pass_2_out;
  wire fifo_cout_drain_PE_7_9_V_full_n_pass_1_out;
  wire fifo_cout_drain_PE_7_9_V_full_n_pass_2_in;
  wire PE_wrapper243_U0_fifo_cout_drain_out_V_write_pass_1_in;
  wire PE_wrapper243_U0_fifo_cout_drain_out_V_write_pass_2_out;
  wire [255:0] PE_wrapper243_U0_fifo_cin_out_V_V_din_pass_1_in;
  wire [255:0] PE_wrapper243_U0_fifo_cin_out_V_V_din_pass_2_out;
  wire fifo_cin_PE_8_9_V_V_full_n_pass_1_out;
  wire fifo_cin_PE_8_9_V_V_full_n_pass_2_in;
  wire PE_wrapper243_U0_fifo_cin_out_V_V_write_pass_1_in;
  wire PE_wrapper243_U0_fifo_cin_out_V_V_write_pass_2_out;
  wire [63:0] cout_drain_IO_L3_out_U0_fifo_cout_drain_out_V_V_din_pass_0_in;
  wire [63:0] cout_drain_IO_L3_out_U0_fifo_cout_drain_out_V_V_din_pass_1_out;
  wire fifo_cout_drain_cout_drain_IO_L3_out_serialize_V_V_full_n_pass_0_out;
  wire fifo_cout_drain_cout_drain_IO_L3_out_serialize_V_V_full_n_pass_1_in;
  wire cout_drain_IO_L3_out_U0_fifo_cout_drain_out_V_V_write_pass_0_in;
  wire cout_drain_IO_L3_out_U0_fifo_cout_drain_out_V_V_write_pass_1_out;
  wire [255:0] PE_wrapper192_U0_fifo_cin_out_V_V_din_pass_0_in;
  wire fifo_cin_PE_4_6_V_V_full_n_pass_0_out;
  wire PE_wrapper192_U0_fifo_cin_out_V_V_write_pass_0_in;
  wire [63:0] cout_drain_IO_L1_out_wrapper471_U0_fifo_cout_drain_out_V_V_din_pass_0_in;
  wire fifo_cout_drain_cout_drain_IO_L1_out_6_7_V_V_full_n_pass_0_out;
  wire cout_drain_IO_L1_out_wrapper471_U0_fifo_cout_drain_out_V_V_write_pass_0_in;
  wire [255:0] PE_wrapper214_U0_fifo_w_out_V_V_din_pass_1_in;
  wire fifo_w_PE_5_5_V_V_full_n_pass_1_out;
  wire PE_wrapper214_U0_fifo_w_out_V_V_write_pass_1_in;
  wire [63:0] cout_drain_IO_L1_out_wrapper490_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_7_4_V_V_full_n_pass_0_in;
  wire cout_drain_IO_L1_out_wrapper490_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper205_U0_fifo_cin_out_V_V_din_pass_0_in;
  wire fifo_cin_PE_5_7_V_V_full_n_pass_0_out;
  wire PE_wrapper205_U0_fifo_cin_out_V_V_write_pass_0_in;
  wire [255:0] PE_wrapper217_U0_fifo_w_out_V_V_din_pass_0_out;
  wire fifo_w_PE_5_8_V_V_full_n_pass_0_in;
  wire PE_wrapper217_U0_fifo_w_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper215_U0_fifo_cin_out_V_V_din_pass_0_out;
  wire fifo_cin_PE_6_5_V_V_full_n_pass_0_in;
  wire PE_wrapper215_U0_fifo_cin_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper227_U0_fifo_w_out_V_V_din_pass_0_in;
  wire fifo_w_PE_6_6_V_V_full_n_pass_0_out;
  wire PE_wrapper227_U0_fifo_w_out_V_V_write_pass_0_in;
  wire [255:0] PE_wrapper228_U0_fifo_cin_out_V_V_din_pass_0_out;
  wire fifo_cin_PE_7_6_V_V_full_n_pass_0_in;
  wire PE_wrapper228_U0_fifo_cin_out_V_V_write_pass_0_out;
  wire [63:0] cout_drain_IO_L1_out_wrapper474_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_6_4_V_V_full_n_pass_0_in;
  wire cout_drain_IO_L1_out_wrapper474_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  wire [63:0] cout_drain_IO_L1_out_wrapper458_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_5_4_V_V_full_n_pass_0_in;
  wire cout_drain_IO_L1_out_wrapper458_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper229_U0_fifo_w_out_V_V_din_pass_0_out;
  wire fifo_w_PE_6_8_V_V_full_n_pass_0_in;
  wire PE_wrapper229_U0_fifo_w_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper202_U0_fifo_w_out_V_V_din_pass_1_in;
  wire fifo_w_PE_4_5_V_V_full_n_pass_1_out;
  wire PE_wrapper202_U0_fifo_w_out_V_V_write_pass_1_in;
  wire [63:0] cout_drain_IO_L1_out_wrapper456_U0_fifo_cout_drain_out_V_V_din_pass_0_in;
  wire fifo_cout_drain_cout_drain_IO_L1_out_5_6_V_V_full_n_pass_0_out;
  wire cout_drain_IO_L1_out_wrapper456_U0_fifo_cout_drain_out_V_V_write_pass_0_in;
  wire [255:0] PE_wrapper229_U0_fifo_cin_out_V_V_din_pass_0_out;
  wire fifo_cin_PE_7_7_V_V_full_n_pass_0_in;
  wire PE_wrapper229_U0_fifo_cin_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper191_U0_fifo_cin_out_V_V_din_pass_0_in;
  wire fifo_cin_PE_4_5_V_V_full_n_pass_0_out;
  wire PE_wrapper191_U0_fifo_cin_out_V_V_write_pass_0_in;
  wire [31:0] PE_wrapper205_U0_fifo_cout_drain_out_V_din_pass_0_in;
  wire fifo_cout_drain_PE_4_7_V_full_n_pass_0_out;
  wire PE_wrapper205_U0_fifo_cout_drain_out_V_write_pass_0_in;
  wire [255:0] PE_wrapper204_U0_fifo_w_out_V_V_din_pass_0_out;
  wire fifo_w_PE_4_7_V_V_full_n_pass_0_in;
  wire PE_wrapper204_U0_fifo_w_out_V_V_write_pass_0_out;
  wire [63:0] cout_drain_IO_L1_out_wrapper487_U0_fifo_cout_drain_out_V_V_din_pass_0_in;
  wire fifo_cout_drain_cout_drain_IO_L1_out_7_7_V_V_full_n_pass_0_out;
  wire cout_drain_IO_L1_out_wrapper487_U0_fifo_cout_drain_out_V_V_write_pass_0_in;
  wire ap_start_Boundary_X4Y8_To_X6Y8_in;
  wire ap_rst_n_Boundary_X4Y8_To_X6Y8_in;
  wire ap_done_Boundary_X4Y8_To_X6Y8_out;
  wire ap_start_Boundary_X4Y10_To_X6Y10_out;
  wire ap_rst_n_Boundary_X4Y10_To_X6Y10_out;
  wire ap_done_Boundary_X4Y10_To_X6Y10_in;
  wire [63:0] kernel0_entry12_U0_cout_V_out_din_pass_4_in;
  wire [63:0] kernel0_entry12_U0_cout_V_out_din_pass_5_out;
  wire cout_V_c_full_n_pass_4_out;
  wire cout_V_c_full_n_pass_5_in;
  wire kernel0_entry12_U0_cout_V_out_write_pass_4_in;
  wire kernel0_entry12_U0_cout_V_out_write_pass_5_out;
  wire [255:0] PE_wrapper243_U0_fifo_w_out_V_V_din_pass_2_in;
  wire [255:0] PE_wrapper243_U0_fifo_w_out_V_V_din_pass_3_out;
  wire fifo_w_PE_7_10_V_V_full_n_pass_2_out;
  wire fifo_w_PE_7_10_V_V_full_n_pass_3_in;
  wire PE_wrapper243_U0_fifo_w_out_V_V_write_pass_2_in;
  wire PE_wrapper243_U0_fifo_w_out_V_V_write_pass_3_out;
  wire [31:0] PE_wrapper243_U0_fifo_cout_drain_out_V_din_pass_2_in;
  wire [31:0] PE_wrapper243_U0_fifo_cout_drain_out_V_din_pass_3_out;
  wire fifo_cout_drain_PE_7_9_V_full_n_pass_2_out;
  wire fifo_cout_drain_PE_7_9_V_full_n_pass_3_in;
  wire PE_wrapper243_U0_fifo_cout_drain_out_V_write_pass_2_in;
  wire PE_wrapper243_U0_fifo_cout_drain_out_V_write_pass_3_out;
  wire [255:0] PE_wrapper243_U0_fifo_cin_out_V_V_din_pass_2_in;
  wire [255:0] PE_wrapper243_U0_fifo_cin_out_V_V_din_pass_3_out;
  wire fifo_cin_PE_8_9_V_V_full_n_pass_2_out;
  wire fifo_cin_PE_8_9_V_V_full_n_pass_3_in;
  wire PE_wrapper243_U0_fifo_cin_out_V_V_write_pass_2_in;
  wire PE_wrapper243_U0_fifo_cin_out_V_V_write_pass_3_out;
  wire [255:0] PE_wrapper182_U0_fifo_w_out_V_V_din_pass_0_in;
  wire [255:0] PE_wrapper182_U0_fifo_w_out_V_V_din_pass_1_out;
  wire fifo_w_PE_2_9_V_V_full_n_pass_0_out;
  wire fifo_w_PE_2_9_V_V_full_n_pass_1_in;
  wire PE_wrapper182_U0_fifo_w_out_V_V_write_pass_0_in;
  wire PE_wrapper182_U0_fifo_w_out_V_V_write_pass_1_out;
  wire [63:0] cout_drain_IO_L3_out_U0_fifo_cout_drain_out_V_V_din_pass_1_in;
  wire [63:0] cout_drain_IO_L3_out_U0_fifo_cout_drain_out_V_V_din_pass_2_out;
  wire fifo_cout_drain_cout_drain_IO_L3_out_serialize_V_V_full_n_pass_1_out;
  wire fifo_cout_drain_cout_drain_IO_L3_out_serialize_V_V_full_n_pass_2_in;
  wire cout_drain_IO_L3_out_U0_fifo_cout_drain_out_V_V_write_pass_1_in;
  wire cout_drain_IO_L3_out_U0_fifo_cout_drain_out_V_V_write_pass_2_out;
  wire [255:0] PE_wrapper194_U0_fifo_w_out_V_V_din_pass_0_in;
  wire [255:0] PE_wrapper194_U0_fifo_w_out_V_V_din_pass_1_out;
  wire fifo_w_PE_3_9_V_V_full_n_pass_0_out;
  wire fifo_w_PE_3_9_V_V_full_n_pass_1_in;
  wire PE_wrapper194_U0_fifo_w_out_V_V_write_pass_0_in;
  wire PE_wrapper194_U0_fifo_w_out_V_V_write_pass_1_out;
  wire [255:0] PE_wrapper253_U0_fifo_cin_out_V_V_din_pass_0_out;
  wire fifo_cin_PE_9_7_V_V_full_n_pass_0_in;
  wire PE_wrapper253_U0_fifo_cin_out_V_V_write_pass_0_out;
  wire [63:0] cout_drain_IO_L1_out_wrapper471_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_6_7_V_V_full_n_pass_0_in;
  wire cout_drain_IO_L1_out_wrapper471_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  wire [31:0] PE_wrapper218_U0_fifo_cout_drain_out_V_din_pass_0_in;
  wire fifo_cout_drain_PE_5_8_V_full_n_pass_0_out;
  wire PE_wrapper218_U0_fifo_cout_drain_out_V_write_pass_0_in;
  wire [255:0] PE_wrapper242_U0_fifo_w_out_V_V_din_pass_0_out;
  wire fifo_w_PE_7_9_V_V_full_n_pass_0_in;
  wire PE_wrapper242_U0_fifo_w_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper230_U0_fifo_w_out_V_V_din_pass_0_out;
  wire fifo_w_PE_6_9_V_V_full_n_pass_0_in;
  wire PE_wrapper230_U0_fifo_w_out_V_V_write_pass_0_out;
  wire [63:0] cout_drain_IO_L1_out_wrapper506_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_8_4_V_V_full_n_pass_0_in;
  wire cout_drain_IO_L1_out_wrapper506_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper252_U0_fifo_cin_out_V_V_din_pass_0_out;
  wire fifo_cin_PE_9_6_V_V_full_n_pass_0_in;
  wire PE_wrapper252_U0_fifo_cin_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper228_U0_fifo_cin_out_V_V_din_pass_0_in;
  wire fifo_cin_PE_7_6_V_V_full_n_pass_0_out;
  wire PE_wrapper228_U0_fifo_cin_out_V_V_write_pass_0_in;
  wire [255:0] PE_wrapper254_U0_fifo_w_out_V_V_din_pass_0_out;
  wire fifo_w_PE_8_9_V_V_full_n_pass_0_in;
  wire PE_wrapper254_U0_fifo_w_out_V_V_write_pass_0_out;
  wire [63:0] cout_drain_IO_L1_out_wrapper501_U0_fifo_cout_drain_out_V_V_din_pass_0_in;
  wire fifo_cout_drain_cout_drain_IO_L1_out_8_9_V_V_full_n_pass_0_out;
  wire cout_drain_IO_L1_out_wrapper501_U0_fifo_cout_drain_out_V_V_write_pass_0_in;
  wire [255:0] PE_wrapper229_U0_fifo_w_out_V_V_din_pass_0_in;
  wire fifo_w_PE_6_8_V_V_full_n_pass_0_out;
  wire PE_wrapper229_U0_fifo_w_out_V_V_write_pass_0_in;
  wire [255:0] PE_wrapper229_U0_fifo_cin_out_V_V_din_pass_0_in;
  wire fifo_cin_PE_7_7_V_V_full_n_pass_0_out;
  wire PE_wrapper229_U0_fifo_cin_out_V_V_write_pass_0_in;
  wire [255:0] PE_wrapper251_U0_fifo_w_out_V_V_din_pass_1_in;
  wire fifo_w_PE_8_6_V_V_full_n_pass_1_out;
  wire PE_wrapper251_U0_fifo_w_out_V_V_write_pass_1_in;
  wire [63:0] cout_drain_IO_L1_out_wrapper485_U0_fifo_cout_drain_out_V_V_din_pass_0_in;
  wire fifo_cout_drain_cout_drain_IO_L1_out_7_9_V_V_full_n_pass_0_out;
  wire cout_drain_IO_L1_out_wrapper485_U0_fifo_cout_drain_out_V_V_write_pass_0_in;
  wire [63:0] cout_drain_IO_L1_out_wrapper487_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_7_7_V_V_full_n_pass_0_in;
  wire cout_drain_IO_L1_out_wrapper487_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  wire [31:0] PE_wrapper206_U0_fifo_cout_drain_out_V_din_pass_0_in;
  wire fifo_cout_drain_PE_4_8_V_full_n_pass_0_out;
  wire PE_wrapper206_U0_fifo_cout_drain_out_V_write_pass_0_in;
  wire [255:0] PE_wrapper218_U0_fifo_cin_out_V_V_din_pass_0_in;
  wire fifo_cin_PE_6_8_V_V_full_n_pass_0_out;
  wire PE_wrapper218_U0_fifo_cin_out_V_V_write_pass_0_in;
  wire [255:0] PE_wrapper239_U0_fifo_w_out_V_V_din_pass_1_in;
  wire fifo_w_PE_7_6_V_V_full_n_pass_1_out;
  wire PE_wrapper239_U0_fifo_w_out_V_V_write_pass_1_in;
  wire [255:0] PE_wrapper254_U0_fifo_cin_out_V_V_din_pass_0_out;
  wire fifo_cin_PE_9_8_V_V_full_n_pass_0_in;
  wire PE_wrapper254_U0_fifo_cin_out_V_V_write_pass_0_out;
  wire [63:0] cout_drain_IO_L1_out_wrapper469_U0_fifo_cout_drain_out_V_V_din_pass_1_in;
  wire fifo_cout_drain_cout_drain_IO_L1_out_6_9_V_V_full_n_pass_1_out;
  wire cout_drain_IO_L1_out_wrapper469_U0_fifo_cout_drain_out_V_V_write_pass_1_in;
  wire ap_start_Boundary_X4Y10_To_X6Y10_in;
  wire ap_rst_n_Boundary_X4Y10_To_X6Y10_in;
  wire ap_done_Boundary_X4Y10_To_X6Y10_out;
  wire ap_start_Boundary_X4Y12_To_X6Y12_out;
  wire ap_rst_n_Boundary_X4Y12_To_X6Y12_out;
  wire ap_done_Boundary_X4Y12_To_X6Y12_in;
  wire [255:0] PE_wrapper242_U0_fifo_w_out_V_V_din_pass_1_in;
  wire [255:0] PE_wrapper242_U0_fifo_w_out_V_V_din_pass_2_out;
  wire fifo_w_PE_7_9_V_V_full_n_pass_1_out;
  wire fifo_w_PE_7_9_V_V_full_n_pass_2_in;
  wire PE_wrapper242_U0_fifo_w_out_V_V_write_pass_1_in;
  wire PE_wrapper242_U0_fifo_w_out_V_V_write_pass_2_out;
  wire [63:0] cout_drain_IO_L1_out_wrapper474_U0_fifo_cout_drain_out_V_V_din_pass_0_in;
  wire [63:0] cout_drain_IO_L1_out_wrapper474_U0_fifo_cout_drain_out_V_V_din_pass_1_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_6_4_V_V_full_n_pass_0_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_6_4_V_V_full_n_pass_1_in;
  wire cout_drain_IO_L1_out_wrapper474_U0_fifo_cout_drain_out_V_V_write_pass_0_in;
  wire cout_drain_IO_L1_out_wrapper474_U0_fifo_cout_drain_out_V_V_write_pass_1_out;
  wire [63:0] cout_drain_IO_L1_out_wrapper458_U0_fifo_cout_drain_out_V_V_din_pass_0_in;
  wire [63:0] cout_drain_IO_L1_out_wrapper458_U0_fifo_cout_drain_out_V_V_din_pass_1_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_5_4_V_V_full_n_pass_0_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_5_4_V_V_full_n_pass_1_in;
  wire cout_drain_IO_L1_out_wrapper458_U0_fifo_cout_drain_out_V_V_write_pass_0_in;
  wire cout_drain_IO_L1_out_wrapper458_U0_fifo_cout_drain_out_V_V_write_pass_1_out;
  wire [255:0] PE_wrapper231_U0_fifo_cin_out_V_V_din_pass_3_in;
  wire [255:0] PE_wrapper231_U0_fifo_cin_out_V_V_din_pass_4_out;
  wire fifo_cin_PE_7_9_V_V_full_n_pass_3_out;
  wire fifo_cin_PE_7_9_V_V_full_n_pass_4_in;
  wire PE_wrapper231_U0_fifo_cin_out_V_V_write_pass_3_in;
  wire PE_wrapper231_U0_fifo_cin_out_V_V_write_pass_4_out;
  wire [255:0] PE_wrapper217_U0_fifo_w_out_V_V_din_pass_0_in;
  wire [255:0] PE_wrapper217_U0_fifo_w_out_V_V_din_pass_1_out;
  wire fifo_w_PE_5_8_V_V_full_n_pass_0_out;
  wire fifo_w_PE_5_8_V_V_full_n_pass_1_in;
  wire PE_wrapper217_U0_fifo_w_out_V_V_write_pass_0_in;
  wire PE_wrapper217_U0_fifo_w_out_V_V_write_pass_1_out;
  wire [255:0] PE_wrapper168_U0_fifo_w_out_V_V_din_pass_0_in;
  wire fifo_w_PE_1_7_V_V_full_n_pass_0_out;
  wire PE_wrapper168_U0_fifo_w_out_V_V_write_pass_0_in;
  wire [255:0] PE_wrapper193_U0_fifo_w_out_V_V_din_pass_0_out;
  wire fifo_w_PE_3_8_V_V_full_n_pass_0_in;
  wire PE_wrapper193_U0_fifo_w_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper181_U0_fifo_w_out_V_V_din_pass_0_out;
  wire fifo_w_PE_2_8_V_V_full_n_pass_0_in;
  wire PE_wrapper181_U0_fifo_w_out_V_V_write_pass_0_out;
  wire [63:0] cout_drain_IO_L2_out561_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  wire fifo_cout_drain_cout_drain_IO_L2_out_7_V_V_full_n_pass_0_in;
  wire cout_drain_IO_L2_out561_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper169_U0_fifo_w_out_V_V_din_pass_0_out;
  wire fifo_w_PE_1_8_V_V_full_n_pass_0_in;
  wire PE_wrapper169_U0_fifo_w_out_V_V_write_pass_0_out;
  wire [255:0] cin_IO_L2_in130_U0_fifo_cin_out_V_V_din_pass_0_in;
  wire fifo_cin_cin_IO_L2_in_7_V_V_full_n_pass_0_out;
  wire cin_IO_L2_in130_U0_fifo_cin_out_V_V_write_pass_0_in;
  wire [255:0] PE_wrapper205_U0_fifo_cin_out_V_V_din_pass_0_out;
  wire fifo_cin_PE_5_7_V_V_full_n_pass_0_in;
  wire PE_wrapper205_U0_fifo_cin_out_V_V_write_pass_0_out;
  wire [63:0] cout_drain_IO_L1_out_wrapper490_U0_fifo_cout_drain_out_V_V_din_pass_0_in;
  wire fifo_cout_drain_cout_drain_IO_L1_out_7_4_V_V_full_n_pass_0_out;
  wire cout_drain_IO_L1_out_wrapper490_U0_fifo_cout_drain_out_V_V_write_pass_0_in;
  wire [255:0] cin_IO_L2_in131_U0_fifo_cin_out_V_V_din_pass_0_out;
  wire fifo_cin_cin_IO_L2_in_8_V_V_full_n_pass_0_in;
  wire cin_IO_L2_in131_U0_fifo_cin_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper156_U0_fifo_w_out_V_V_din_pass_0_in;
  wire fifo_w_PE_0_7_V_V_full_n_pass_0_out;
  wire PE_wrapper156_U0_fifo_w_out_V_V_write_pass_0_in;
  wire [255:0] PE_wrapper157_U0_fifo_w_out_V_V_din_pass_0_out;
  wire fifo_w_PE_0_8_V_V_full_n_pass_0_in;
  wire PE_wrapper157_U0_fifo_w_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper192_U0_fifo_w_out_V_V_din_pass_1_in;
  wire fifo_w_PE_3_7_V_V_full_n_pass_1_out;
  wire PE_wrapper192_U0_fifo_w_out_V_V_write_pass_1_in;
  wire [63:0] cout_drain_IO_L2_out560_U0_fifo_cout_drain_out_V_V_din_pass_0_in;
  wire fifo_cout_drain_cout_drain_IO_L2_out_8_V_V_full_n_pass_0_out;
  wire cout_drain_IO_L2_out560_U0_fifo_cout_drain_out_V_V_write_pass_0_in;
  wire [63:0] cout_drain_IO_L3_out_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  wire fifo_cout_drain_cout_drain_IO_L3_out_serialize_V_V_full_n_pass_0_in;
  wire cout_drain_IO_L3_out_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper180_U0_fifo_w_out_V_V_din_pass_0_in;
  wire fifo_w_PE_2_7_V_V_full_n_pass_0_out;
  wire PE_wrapper180_U0_fifo_w_out_V_V_write_pass_0_in;
  wire [31:0] PE_wrapper205_U0_fifo_cout_drain_out_V_din_pass_0_out;
  wire fifo_cout_drain_PE_4_7_V_full_n_pass_0_in;
  wire PE_wrapper205_U0_fifo_cout_drain_out_V_write_pass_0_out;
  wire [255:0] PE_wrapper205_U0_fifo_w_out_V_V_din_pass_0_out;
  wire fifo_w_PE_4_8_V_V_full_n_pass_0_in;
  wire PE_wrapper205_U0_fifo_w_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper204_U0_fifo_w_out_V_V_din_pass_0_in;
  wire fifo_w_PE_4_7_V_V_full_n_pass_0_out;
  wire PE_wrapper204_U0_fifo_w_out_V_V_write_pass_0_in;
  wire [63:0] cout_drain_IO_L2_out568_U0_fifo_cout_drain_out_V_V_din_pass_3_in;
  wire fifo_cout_drain_cout_drain_IO_L2_out_0_V_V_full_n_pass_3_out;
  wire cout_drain_IO_L2_out568_U0_fifo_cout_drain_out_V_V_write_pass_3_in;
  wire ap_start_Boundary_X6Y8_To_X8Y8_in;
  wire ap_rst_n_Boundary_X6Y8_To_X8Y8_in;
  wire ap_done_Boundary_X6Y8_To_X8Y8_out;
  wire ap_start_Boundary_X6Y10_To_X8Y10_out;
  wire ap_rst_n_Boundary_X6Y10_To_X8Y10_out;
  wire ap_done_Boundary_X6Y10_To_X8Y10_in;
  wire [255:0] PE_wrapper242_U0_fifo_w_out_V_V_din_pass_0_in;
  wire [255:0] PE_wrapper242_U0_fifo_w_out_V_V_din_pass_1_out;
  wire fifo_w_PE_7_9_V_V_full_n_pass_0_out;
  wire fifo_w_PE_7_9_V_V_full_n_pass_1_in;
  wire PE_wrapper242_U0_fifo_w_out_V_V_write_pass_0_in;
  wire PE_wrapper242_U0_fifo_w_out_V_V_write_pass_1_out;
  wire [255:0] PE_wrapper231_U0_fifo_cin_out_V_V_din_pass_2_in;
  wire [255:0] PE_wrapper231_U0_fifo_cin_out_V_V_din_pass_3_out;
  wire fifo_cin_PE_7_9_V_V_full_n_pass_2_out;
  wire fifo_cin_PE_7_9_V_V_full_n_pass_3_in;
  wire PE_wrapper231_U0_fifo_cin_out_V_V_write_pass_2_in;
  wire PE_wrapper231_U0_fifo_cin_out_V_V_write_pass_3_out;
  wire [255:0] PE_wrapper158_U0_fifo_w_out_V_V_din_pass_0_out;
  wire fifo_w_PE_0_9_V_V_full_n_pass_0_in;
  wire PE_wrapper158_U0_fifo_w_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper193_U0_fifo_w_out_V_V_din_pass_0_in;
  wire fifo_w_PE_3_8_V_V_full_n_pass_0_out;
  wire PE_wrapper193_U0_fifo_w_out_V_V_write_pass_0_in;
  wire [255:0] PE_wrapper170_U0_fifo_w_out_V_V_din_pass_0_out;
  wire fifo_w_PE_1_9_V_V_full_n_pass_0_in;
  wire PE_wrapper170_U0_fifo_w_out_V_V_write_pass_0_out;
  wire [63:0] cout_drain_IO_L2_out559_U0_fifo_cout_drain_out_V_V_din_pass_0_in;
  wire fifo_cout_drain_cout_drain_IO_L2_out_9_V_V_full_n_pass_0_out;
  wire cout_drain_IO_L2_out559_U0_fifo_cout_drain_out_V_V_write_pass_0_in;
  wire [255:0] PE_wrapper181_U0_fifo_w_out_V_V_din_pass_0_in;
  wire fifo_w_PE_2_8_V_V_full_n_pass_0_out;
  wire PE_wrapper181_U0_fifo_w_out_V_V_write_pass_0_in;
  wire [255:0] PE_wrapper206_U0_fifo_w_out_V_V_din_pass_0_out;
  wire fifo_w_PE_4_9_V_V_full_n_pass_0_in;
  wire PE_wrapper206_U0_fifo_w_out_V_V_write_pass_0_out;
  wire [255:0] cin_IO_L2_in132_U0_fifo_cin_out_V_V_din_pass_0_out;
  wire fifo_cin_cin_IO_L2_in_9_V_V_full_n_pass_0_in;
  wire cin_IO_L2_in132_U0_fifo_cin_out_V_V_write_pass_0_out;
  wire [31:0] PE_wrapper218_U0_fifo_cout_drain_out_V_din_pass_0_out;
  wire fifo_cout_drain_PE_5_8_V_full_n_pass_0_in;
  wire PE_wrapper218_U0_fifo_cout_drain_out_V_write_pass_0_out;
  wire [63:0] cout_drain_IO_L1_out_wrapper506_U0_fifo_cout_drain_out_V_V_din_pass_0_in;
  wire fifo_cout_drain_cout_drain_IO_L1_out_8_4_V_V_full_n_pass_0_out;
  wire cout_drain_IO_L1_out_wrapper506_U0_fifo_cout_drain_out_V_V_write_pass_0_in;
  wire [255:0] PE_wrapper169_U0_fifo_w_out_V_V_din_pass_0_in;
  wire fifo_w_PE_1_8_V_V_full_n_pass_0_out;
  wire PE_wrapper169_U0_fifo_w_out_V_V_write_pass_0_in;
  wire [255:0] PE_wrapper217_U0_fifo_w_out_V_V_din_pass_1_in;
  wire fifo_w_PE_5_8_V_V_full_n_pass_1_out;
  wire PE_wrapper217_U0_fifo_w_out_V_V_write_pass_1_in;
  wire [255:0] cin_IO_L2_in131_U0_fifo_cin_out_V_V_din_pass_0_in;
  wire fifo_cin_cin_IO_L2_in_8_V_V_full_n_pass_0_out;
  wire cin_IO_L2_in131_U0_fifo_cin_out_V_V_write_pass_0_in;
  wire [255:0] PE_wrapper157_U0_fifo_w_out_V_V_din_pass_0_in;
  wire fifo_w_PE_0_8_V_V_full_n_pass_0_out;
  wire PE_wrapper157_U0_fifo_w_out_V_V_write_pass_0_in;
  wire [255:0] PE_wrapper182_U0_fifo_w_out_V_V_din_pass_0_out;
  wire fifo_w_PE_2_9_V_V_full_n_pass_0_in;
  wire PE_wrapper182_U0_fifo_w_out_V_V_write_pass_0_out;
  wire [63:0] cout_drain_IO_L2_out560_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  wire fifo_cout_drain_cout_drain_IO_L2_out_8_V_V_full_n_pass_0_in;
  wire cout_drain_IO_L2_out560_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper205_U0_fifo_w_out_V_V_din_pass_0_in;
  wire fifo_w_PE_4_8_V_V_full_n_pass_0_out;
  wire PE_wrapper205_U0_fifo_w_out_V_V_write_pass_0_in;
  wire [255:0] PE_wrapper218_U0_fifo_w_out_V_V_din_pass_0_out;
  wire fifo_w_PE_5_9_V_V_full_n_pass_0_in;
  wire PE_wrapper218_U0_fifo_w_out_V_V_write_pass_0_out;
  wire [31:0] PE_wrapper206_U0_fifo_cout_drain_out_V_din_pass_0_out;
  wire fifo_cout_drain_PE_4_8_V_full_n_pass_0_in;
  wire PE_wrapper206_U0_fifo_cout_drain_out_V_write_pass_0_out;
  wire [255:0] PE_wrapper218_U0_fifo_cin_out_V_V_din_pass_0_out;
  wire fifo_cin_PE_6_8_V_V_full_n_pass_0_in;
  wire PE_wrapper218_U0_fifo_cin_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper194_U0_fifo_w_out_V_V_din_pass_0_out;
  wire fifo_w_PE_3_9_V_V_full_n_pass_0_in;
  wire PE_wrapper194_U0_fifo_w_out_V_V_write_pass_0_out;
  wire ap_start_Boundary_X6Y10_To_X8Y10_in;
  wire ap_rst_n_Boundary_X6Y10_To_X8Y10_in;
  wire ap_done_Boundary_X6Y10_To_X8Y10_out;
  wire ap_start_Boundary_X6Y12_To_X8Y12_out;
  wire ap_rst_n_Boundary_X6Y12_To_X8Y12_out;
  wire ap_done_Boundary_X6Y12_To_X8Y12_in;
  wire [255:0] PE_wrapper256_U0_fifo_cin_out_V_V_din_pass_0_in;
  wire [255:0] PE_wrapper256_U0_fifo_cin_out_V_V_din_pass_1_out;
  wire fifo_cin_PE_9_10_V_V_full_n_pass_0_out;
  wire fifo_cin_PE_9_10_V_V_full_n_pass_1_in;
  wire PE_wrapper256_U0_fifo_cin_out_V_V_write_pass_0_in;
  wire PE_wrapper256_U0_fifo_cin_out_V_V_write_pass_1_out;
  wire [255:0] PE_wrapper257_U0_fifo_cin_out_V_V_din_pass_0_in;
  wire [255:0] PE_wrapper257_U0_fifo_cin_out_V_V_din_pass_1_out;
  wire fifo_cin_PE_9_11_V_V_full_n_pass_0_out;
  wire fifo_cin_PE_9_11_V_V_full_n_pass_1_in;
  wire PE_wrapper257_U0_fifo_cin_out_V_V_write_pass_0_in;
  wire PE_wrapper257_U0_fifo_cin_out_V_V_write_pass_1_out;
  wire [63:0] cout_drain_IO_L1_out_wrapper551_U0_fifo_cout_drain_out_V_V_din_pass_0_in;
  wire [63:0] cout_drain_IO_L1_out_wrapper551_U0_fifo_cout_drain_out_V_V_din_pass_1_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_11_6_V_V_full_n_pass_0_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_11_6_V_V_full_n_pass_1_in;
  wire cout_drain_IO_L1_out_wrapper551_U0_fifo_cout_drain_out_V_V_write_pass_0_in;
  wire cout_drain_IO_L1_out_wrapper551_U0_fifo_cout_drain_out_V_V_write_pass_1_out;
  wire [255:0] PE_wrapper161_U0_fifo_cin_out_V_V_din_pass_0_in;
  wire [255:0] PE_wrapper161_U0_fifo_cin_out_V_V_din_pass_1_out;
  wire fifo_cin_PE_1_11_V_V_full_n_pass_0_out;
  wire fifo_cin_PE_1_11_V_V_full_n_pass_1_in;
  wire PE_wrapper161_U0_fifo_cin_out_V_V_write_pass_0_in;
  wire PE_wrapper161_U0_fifo_cin_out_V_V_write_pass_1_out;
  wire [31:0] PE_wrapper185_U0_fifo_cout_drain_out_V_din_pass_0_in;
  wire [31:0] PE_wrapper185_U0_fifo_cout_drain_out_V_din_pass_1_out;
  wire fifo_cout_drain_PE_2_11_V_full_n_pass_0_out;
  wire fifo_cout_drain_PE_2_11_V_full_n_pass_1_in;
  wire PE_wrapper185_U0_fifo_cout_drain_out_V_write_pass_0_in;
  wire PE_wrapper185_U0_fifo_cout_drain_out_V_write_pass_1_out;
  wire [63:0] cout_drain_IO_L1_out_wrapper518_U0_fifo_cout_drain_out_V_V_din_pass_0_in;
  wire [63:0] cout_drain_IO_L1_out_wrapper518_U0_fifo_cout_drain_out_V_V_din_pass_1_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_9_8_V_V_full_n_pass_0_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_9_8_V_V_full_n_pass_1_in;
  wire cout_drain_IO_L1_out_wrapper518_U0_fifo_cout_drain_out_V_V_write_pass_0_in;
  wire cout_drain_IO_L1_out_wrapper518_U0_fifo_cout_drain_out_V_V_write_pass_1_out;
  wire [63:0] cout_drain_IO_L1_out_wrapper534_U0_fifo_cout_drain_out_V_V_din_pass_0_in;
  wire [63:0] cout_drain_IO_L1_out_wrapper534_U0_fifo_cout_drain_out_V_V_din_pass_1_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_10_8_V_V_full_n_pass_0_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_10_8_V_V_full_n_pass_1_in;
  wire cout_drain_IO_L1_out_wrapper534_U0_fifo_cout_drain_out_V_V_write_pass_0_in;
  wire cout_drain_IO_L1_out_wrapper534_U0_fifo_cout_drain_out_V_V_write_pass_1_out;
  wire [31:0] PE_wrapper197_U0_fifo_cout_drain_out_V_din_pass_0_in;
  wire [31:0] PE_wrapper197_U0_fifo_cout_drain_out_V_din_pass_1_out;
  wire fifo_cout_drain_PE_3_11_V_full_n_pass_0_out;
  wire fifo_cout_drain_PE_3_11_V_full_n_pass_1_in;
  wire PE_wrapper197_U0_fifo_cout_drain_out_V_write_pass_0_in;
  wire PE_wrapper197_U0_fifo_cout_drain_out_V_write_pass_1_out;
  wire [63:0] cout_drain_IO_L1_out_wrapper523_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_9_3_V_V_full_n_pass_0_in;
  wire cout_drain_IO_L1_out_wrapper523_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  wire [63:0] cout_drain_IO_L1_out_wrapper535_U0_fifo_cout_drain_out_V_V_din_pass_0_in;
  wire fifo_cout_drain_cout_drain_IO_L1_out_10_7_V_V_full_n_pass_0_out;
  wire cout_drain_IO_L1_out_wrapper535_U0_fifo_cout_drain_out_V_V_write_pass_0_in;
  wire [63:0] cout_drain_IO_L1_out_wrapper537_U0_fifo_cout_drain_out_V_V_din_pass_0_in;
  wire fifo_cout_drain_cout_drain_IO_L1_out_10_5_V_V_full_n_pass_0_out;
  wire cout_drain_IO_L1_out_wrapper537_U0_fifo_cout_drain_out_V_V_write_pass_0_in;
  wire [63:0] cout_drain_IO_L1_out_wrapper555_U0_fifo_cout_drain_out_V_V_din_pass_0_in;
  wire fifo_cout_drain_cout_drain_IO_L1_out_11_2_V_V_full_n_pass_0_out;
  wire cout_drain_IO_L1_out_wrapper555_U0_fifo_cout_drain_out_V_V_write_pass_0_in;
  wire [255:0] PE_wrapper196_U0_fifo_cin_out_V_V_din_pass_0_out;
  wire fifo_cin_PE_4_10_V_V_full_n_pass_0_in;
  wire PE_wrapper196_U0_fifo_cin_out_V_V_write_pass_0_out;
  wire [63:0] cout_drain_IO_L1_out_wrapper556_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_11_1_V_V_full_n_pass_0_in;
  wire cout_drain_IO_L1_out_wrapper556_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  wire [63:0] cout_drain_IO_L1_out_wrapper539_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_10_3_V_V_full_n_pass_0_in;
  wire cout_drain_IO_L1_out_wrapper539_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper231_U0_fifo_w_out_V_V_din_pass_0_out;
  wire fifo_w_PE_6_10_V_V_full_n_pass_0_in;
  wire PE_wrapper231_U0_fifo_w_out_V_V_write_pass_0_out;
  wire [31:0] PE_wrapper231_U0_fifo_cout_drain_out_V_din_pass_0_out;
  wire fifo_cout_drain_PE_6_9_V_full_n_pass_0_in;
  wire PE_wrapper231_U0_fifo_cout_drain_out_V_write_pass_0_out;
  wire [255:0] PE_wrapper230_U0_fifo_w_out_V_V_din_pass_1_in;
  wire fifo_w_PE_6_9_V_V_full_n_pass_1_out;
  wire PE_wrapper230_U0_fifo_w_out_V_V_write_pass_1_in;
  wire [63:0] cout_drain_IO_L2_out558_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  wire fifo_cout_drain_cout_drain_IO_L2_out_10_V_V_full_n_pass_0_in;
  wire cout_drain_IO_L2_out558_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  wire [31:0] PE_wrapper221_U0_fifo_cout_drain_out_V_din_pass_0_out;
  wire fifo_cout_drain_PE_5_11_V_full_n_pass_0_in;
  wire PE_wrapper221_U0_fifo_cout_drain_out_V_write_pass_0_out;
  wire [255:0] PE_wrapper184_U0_fifo_w_out_V_V_din_pass_0_out;
  wire fifo_w_PE_2_11_V_V_full_n_pass_0_in;
  wire PE_wrapper184_U0_fifo_w_out_V_V_write_pass_0_out;
  wire [31:0] PE_wrapper232_U0_fifo_cout_drain_out_V_din_pass_0_in;
  wire fifo_cout_drain_PE_6_10_V_full_n_pass_0_out;
  wire PE_wrapper232_U0_fifo_cout_drain_out_V_write_pass_0_in;
  wire [63:0] cout_drain_IO_L1_out_wrapper522_U0_fifo_cout_drain_out_V_V_din_pass_1_in;
  wire fifo_cout_drain_cout_drain_IO_L1_out_9_4_V_V_full_n_pass_1_out;
  wire cout_drain_IO_L1_out_wrapper522_U0_fifo_cout_drain_out_V_V_write_pass_1_in;
  wire [255:0] PE_wrapper196_U0_fifo_w_out_V_V_din_pass_0_out;
  wire fifo_w_PE_3_11_V_V_full_n_pass_0_in;
  wire PE_wrapper196_U0_fifo_w_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper209_U0_fifo_w_out_V_V_din_pass_0_out;
  wire fifo_w_PE_4_12_V_V_full_n_pass_0_in;
  wire PE_wrapper209_U0_fifo_w_out_V_V_write_pass_0_out;
  wire [63:0] cout_drain_IO_L1_out_wrapper552_U0_fifo_cout_drain_out_V_V_din_pass_0_in;
  wire fifo_cout_drain_cout_drain_IO_L1_out_11_5_V_V_full_n_pass_0_out;
  wire cout_drain_IO_L1_out_wrapper552_U0_fifo_cout_drain_out_V_V_write_pass_0_in;
  wire [255:0] PE_wrapper233_U0_fifo_cin_out_V_V_din_pass_0_out;
  wire fifo_cin_PE_7_11_V_V_full_n_pass_0_in;
  wire PE_wrapper233_U0_fifo_cin_out_V_V_write_pass_0_out;
  wire [31:0] PE_wrapper184_U0_fifo_cout_drain_out_V_din_pass_0_out;
  wire fifo_cout_drain_PE_2_10_V_full_n_pass_0_in;
  wire PE_wrapper184_U0_fifo_cout_drain_out_V_write_pass_0_out;
  wire [63:0] cout_drain_IO_L2_out_boundary_U0_fifo_cout_drain_out_V_V_din_pass_0_in;
  wire fifo_cout_drain_cout_drain_IO_L2_out_11_V_V_full_n_pass_0_out;
  wire cout_drain_IO_L2_out_boundary_U0_fifo_cout_drain_out_V_V_write_pass_0_in;
  wire [255:0] PE_wrapper197_U0_fifo_cin_out_V_V_din_pass_0_in;
  wire fifo_cin_PE_4_11_V_V_full_n_pass_0_out;
  wire PE_wrapper197_U0_fifo_cin_out_V_V_write_pass_0_in;
  wire [63:0] cout_drain_IO_L1_out_wrapper542_U0_fifo_cout_drain_out_V_V_din_pass_1_in;
  wire fifo_cout_drain_cout_drain_IO_L1_out_10_0_V_V_full_n_pass_1_out;
  wire cout_drain_IO_L1_out_wrapper542_U0_fifo_cout_drain_out_V_V_write_pass_1_in;
  wire [255:0] PE_wrapper219_U0_fifo_cin_out_V_V_din_pass_1_in;
  wire fifo_cin_PE_6_9_V_V_full_n_pass_1_out;
  wire PE_wrapper219_U0_fifo_cin_out_V_V_write_pass_1_in;
  wire [31:0] PE_wrapper173_U0_fifo_cout_drain_out_V_din_pass_0_in;
  wire fifo_cout_drain_PE_1_11_V_full_n_pass_0_out;
  wire PE_wrapper173_U0_fifo_cout_drain_out_V_write_pass_0_in;
  wire [63:0] cout_drain_IO_L1_out_wrapper549_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_11_8_V_V_full_n_pass_0_in;
  wire cout_drain_IO_L1_out_wrapper549_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper172_U0_fifo_cin_out_V_V_din_pass_1_in;
  wire fifo_cin_PE_2_10_V_V_full_n_pass_1_out;
  wire PE_wrapper172_U0_fifo_cin_out_V_V_write_pass_1_in;
  wire [255:0] PE_wrapper195_U0_fifo_cin_out_V_V_din_pass_0_out;
  wire fifo_cin_PE_4_9_V_V_full_n_pass_0_in;
  wire PE_wrapper195_U0_fifo_cin_out_V_V_write_pass_0_out;
  wire [63:0] cout_drain_IO_L1_out_wrapper536_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_10_6_V_V_full_n_pass_0_in;
  wire cout_drain_IO_L1_out_wrapper536_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  wire [31:0] PE_wrapper208_U0_fifo_cout_drain_out_V_din_pass_0_in;
  wire fifo_cout_drain_PE_4_10_V_full_n_pass_0_out;
  wire PE_wrapper208_U0_fifo_cout_drain_out_V_write_pass_0_in;
  wire [255:0] PE_wrapper220_U0_fifo_w_out_V_V_din_pass_0_in;
  wire fifo_w_PE_5_11_V_V_full_n_pass_0_out;
  wire PE_wrapper220_U0_fifo_w_out_V_V_write_pass_0_in;
  wire [255:0] cin_IO_L2_in134_U0_fifo_cin_out_V_V_din_pass_1_in;
  wire fifo_cin_cin_IO_L2_in_11_V_V_full_n_pass_1_out;
  wire cin_IO_L2_in134_U0_fifo_cin_out_V_V_write_pass_1_in;
  wire [63:0] cout_drain_IO_L1_out_wrapper520_U0_fifo_cout_drain_out_V_V_din_pass_0_in;
  wire fifo_cout_drain_cout_drain_IO_L1_out_9_6_V_V_full_n_pass_0_out;
  wire cout_drain_IO_L1_out_wrapper520_U0_fifo_cout_drain_out_V_V_write_pass_0_in;
  wire [31:0] PE_wrapper257_U0_fifo_cout_drain_out_V_din_pass_0_in;
  wire fifo_cout_drain_PE_8_11_V_full_n_pass_0_out;
  wire PE_wrapper257_U0_fifo_cout_drain_out_V_write_pass_0_in;
  wire [255:0] cin_IO_L2_in_boundary_U0_fifo_cin_local_out_V_V_din_pass_0_out;
  wire fifo_cin_PE_0_11_V_V_full_n_pass_0_in;
  wire cin_IO_L2_in_boundary_U0_fifo_cin_local_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper232_U0_fifo_w_out_V_V_din_pass_0_in;
  wire fifo_w_PE_6_11_V_V_full_n_pass_0_out;
  wire PE_wrapper232_U0_fifo_w_out_V_V_write_pass_0_in;
  wire [255:0] PE_wrapper183_U0_fifo_w_out_V_V_din_pass_0_in;
  wire fifo_w_PE_2_10_V_V_full_n_pass_0_out;
  wire PE_wrapper183_U0_fifo_w_out_V_V_write_pass_0_in;
  wire [255:0] PE_wrapper221_U0_fifo_w_out_V_V_din_pass_0_out;
  wire fifo_w_PE_5_12_V_V_full_n_pass_0_in;
  wire PE_wrapper221_U0_fifo_w_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper208_U0_fifo_w_out_V_V_din_pass_0_in;
  wire fifo_w_PE_4_11_V_V_full_n_pass_0_out;
  wire PE_wrapper208_U0_fifo_w_out_V_V_write_pass_0_in;
  wire [31:0] PE_wrapper233_U0_fifo_cout_drain_out_V_din_pass_0_out;
  wire fifo_cout_drain_PE_6_11_V_full_n_pass_0_in;
  wire PE_wrapper233_U0_fifo_cout_drain_out_V_write_pass_0_out;
  wire [255:0] PE_wrapper183_U0_fifo_cin_out_V_V_din_pass_0_in;
  wire fifo_cin_PE_3_9_V_V_full_n_pass_0_out;
  wire PE_wrapper183_U0_fifo_cin_out_V_V_write_pass_0_in;
  wire [255:0] PE_wrapper194_U0_fifo_w_out_V_V_din_pass_2_in;
  wire fifo_w_PE_3_9_V_V_full_n_pass_2_out;
  wire PE_wrapper194_U0_fifo_w_out_V_V_write_pass_2_in;
  wire [255:0] PE_wrapper231_U0_fifo_cin_out_V_V_din_pass_0_out;
  wire fifo_cin_PE_7_9_V_V_full_n_pass_0_in;
  wire PE_wrapper231_U0_fifo_cin_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper185_U0_fifo_w_out_V_V_din_pass_0_in;
  wire fifo_w_PE_2_12_V_V_full_n_pass_0_out;
  wire PE_wrapper185_U0_fifo_w_out_V_V_write_pass_0_in;
  wire [63:0] cout_drain_IO_L1_out_wrapper548_U0_fifo_cout_drain_out_V_V_din_pass_1_in;
  wire fifo_cout_drain_cout_drain_IO_L1_out_11_9_V_V_full_n_pass_1_out;
  wire cout_drain_IO_L1_out_wrapper548_U0_fifo_cout_drain_out_V_V_write_pass_1_in;
  wire [63:0] cout_drain_IO_L1_out_wrapper521_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_9_5_V_V_full_n_pass_0_in;
  wire cout_drain_IO_L1_out_wrapper521_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  wire [31:0] PE_wrapper219_U0_fifo_cout_drain_out_V_din_pass_1_in;
  wire fifo_cout_drain_PE_5_9_V_full_n_pass_1_out;
  wire PE_wrapper219_U0_fifo_cout_drain_out_V_write_pass_1_in;
  wire [63:0] cout_drain_IO_L1_out_wrapper553_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_11_4_V_V_full_n_pass_0_in;
  wire cout_drain_IO_L1_out_wrapper553_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  wire ap_start_Boundary_X4Y14_To_X6Y14_in;
  wire ap_rst_n_Boundary_X4Y14_To_X6Y14_in;
  wire ap_done_Boundary_X4Y14_To_X6Y14_out;
  wire [255:0] PE_wrapper231_U0_fifo_cin_out_V_V_din_pass_1_in;
  wire [255:0] PE_wrapper231_U0_fifo_cin_out_V_V_din_pass_2_out;
  wire fifo_cin_PE_7_9_V_V_full_n_pass_1_out;
  wire fifo_cin_PE_7_9_V_V_full_n_pass_2_in;
  wire PE_wrapper231_U0_fifo_cin_out_V_V_write_pass_1_in;
  wire PE_wrapper231_U0_fifo_cin_out_V_V_write_pass_2_out;
  wire [255:0] PE_wrapper244_U0_fifo_cin_out_V_V_din_pass_0_in;
  wire [255:0] PE_wrapper244_U0_fifo_cin_out_V_V_din_pass_1_out;
  wire fifo_cin_PE_8_10_V_V_full_n_pass_0_out;
  wire fifo_cin_PE_8_10_V_V_full_n_pass_1_in;
  wire PE_wrapper244_U0_fifo_cin_out_V_V_write_pass_0_in;
  wire PE_wrapper244_U0_fifo_cin_out_V_V_write_pass_1_out;
  wire [255:0] PE_wrapper173_U0_fifo_w_out_V_V_din_pass_0_in;
  wire [255:0] PE_wrapper173_U0_fifo_w_out_V_V_din_pass_1_out;
  wire fifo_w_PE_1_12_V_V_full_n_pass_0_out;
  wire fifo_w_PE_1_12_V_V_full_n_pass_1_in;
  wire PE_wrapper173_U0_fifo_w_out_V_V_write_pass_0_in;
  wire PE_wrapper173_U0_fifo_w_out_V_V_write_pass_1_out;
  wire [31:0] PE_wrapper255_U0_fifo_cout_drain_out_V_din_pass_0_in;
  wire [31:0] PE_wrapper255_U0_fifo_cout_drain_out_V_din_pass_1_out;
  wire fifo_cout_drain_PE_8_9_V_full_n_pass_0_out;
  wire fifo_cout_drain_PE_8_9_V_full_n_pass_1_in;
  wire PE_wrapper255_U0_fifo_cout_drain_out_V_write_pass_0_in;
  wire PE_wrapper255_U0_fifo_cout_drain_out_V_write_pass_1_out;
  wire [255:0] PE_wrapper244_U0_fifo_w_out_V_V_din_pass_0_in;
  wire [255:0] PE_wrapper244_U0_fifo_w_out_V_V_din_pass_1_out;
  wire fifo_w_PE_7_11_V_V_full_n_pass_0_out;
  wire fifo_w_PE_7_11_V_V_full_n_pass_1_in;
  wire PE_wrapper244_U0_fifo_w_out_V_V_write_pass_0_in;
  wire PE_wrapper244_U0_fifo_w_out_V_V_write_pass_1_out;
  wire [63:0] cout_drain_IO_L1_out_wrapper517_U0_fifo_cout_drain_out_V_V_din_pass_1_in;
  wire [63:0] cout_drain_IO_L1_out_wrapper517_U0_fifo_cout_drain_out_V_V_din_pass_2_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_9_9_V_V_full_n_pass_1_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_9_9_V_V_full_n_pass_2_in;
  wire cout_drain_IO_L1_out_wrapper517_U0_fifo_cout_drain_out_V_V_write_pass_1_in;
  wire cout_drain_IO_L1_out_wrapper517_U0_fifo_cout_drain_out_V_V_write_pass_2_out;
  wire [255:0] PE_wrapper255_U0_fifo_w_out_V_V_din_pass_0_in;
  wire [255:0] PE_wrapper255_U0_fifo_w_out_V_V_din_pass_1_out;
  wire fifo_w_PE_8_10_V_V_full_n_pass_0_out;
  wire fifo_w_PE_8_10_V_V_full_n_pass_1_in;
  wire PE_wrapper255_U0_fifo_w_out_V_V_write_pass_0_in;
  wire PE_wrapper255_U0_fifo_w_out_V_V_write_pass_1_out;
  wire [255:0] PE_wrapper173_U0_fifo_cin_out_V_V_din_pass_0_in;
  wire [255:0] PE_wrapper173_U0_fifo_cin_out_V_V_din_pass_1_out;
  wire fifo_cin_PE_2_11_V_V_full_n_pass_0_out;
  wire fifo_cin_PE_2_11_V_V_full_n_pass_1_in;
  wire PE_wrapper173_U0_fifo_cin_out_V_V_write_pass_0_in;
  wire PE_wrapper173_U0_fifo_cin_out_V_V_write_pass_1_out;
  wire [63:0] cout_drain_IO_L1_out_wrapper533_U0_fifo_cout_drain_out_V_V_din_pass_1_in;
  wire [63:0] cout_drain_IO_L1_out_wrapper533_U0_fifo_cout_drain_out_V_V_din_pass_2_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_10_9_V_V_full_n_pass_1_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_10_9_V_V_full_n_pass_2_in;
  wire cout_drain_IO_L1_out_wrapper533_U0_fifo_cout_drain_out_V_V_write_pass_1_in;
  wire cout_drain_IO_L1_out_wrapper533_U0_fifo_cout_drain_out_V_V_write_pass_2_out;
  wire [255:0] PE_wrapper158_U0_fifo_w_out_V_V_din_pass_0_in;
  wire fifo_w_PE_0_9_V_V_full_n_pass_0_out;
  wire PE_wrapper158_U0_fifo_w_out_V_V_write_pass_0_in;
  wire [63:0] cout_drain_IO_L1_out_wrapper523_U0_fifo_cout_drain_out_V_V_din_pass_1_in;
  wire fifo_cout_drain_cout_drain_IO_L1_out_9_3_V_V_full_n_pass_1_out;
  wire cout_drain_IO_L1_out_wrapper523_U0_fifo_cout_drain_out_V_V_write_pass_1_in;
  wire [255:0] PE_wrapper219_U0_fifo_w_out_V_V_din_pass_0_out;
  wire fifo_w_PE_5_10_V_V_full_n_pass_0_in;
  wire PE_wrapper219_U0_fifo_w_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper170_U0_fifo_w_out_V_V_din_pass_0_in;
  wire fifo_w_PE_1_9_V_V_full_n_pass_0_out;
  wire PE_wrapper170_U0_fifo_w_out_V_V_write_pass_0_in;
  wire [255:0] PE_wrapper171_U0_fifo_cin_out_V_V_din_pass_0_out;
  wire fifo_cin_PE_2_9_V_V_full_n_pass_0_in;
  wire PE_wrapper171_U0_fifo_cin_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper172_U0_fifo_w_out_V_V_din_pass_0_out;
  wire fifo_w_PE_1_11_V_V_full_n_pass_0_in;
  wire PE_wrapper172_U0_fifo_w_out_V_V_write_pass_0_out;
  wire [63:0] cout_drain_IO_L2_out559_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  wire fifo_cout_drain_cout_drain_IO_L2_out_9_V_V_full_n_pass_0_in;
  wire cout_drain_IO_L2_out559_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper206_U0_fifo_w_out_V_V_din_pass_0_in;
  wire fifo_w_PE_4_9_V_V_full_n_pass_0_out;
  wire PE_wrapper206_U0_fifo_w_out_V_V_write_pass_0_in;
  wire [255:0] cin_IO_L2_in132_U0_fifo_cin_out_V_V_din_pass_0_in;
  wire fifo_cin_cin_IO_L2_in_9_V_V_full_n_pass_0_out;
  wire cin_IO_L2_in132_U0_fifo_cin_out_V_V_write_pass_0_in;
  wire [255:0] PE_wrapper160_U0_fifo_w_out_V_V_din_pass_0_out;
  wire fifo_w_PE_0_11_V_V_full_n_pass_0_in;
  wire PE_wrapper160_U0_fifo_w_out_V_V_write_pass_0_out;
  wire [63:0] cout_drain_IO_L2_out558_U0_fifo_cout_drain_out_V_V_din_pass_1_in;
  wire fifo_cout_drain_cout_drain_IO_L2_out_10_V_V_full_n_pass_1_out;
  wire cout_drain_IO_L2_out558_U0_fifo_cout_drain_out_V_V_write_pass_1_in;
  wire [255:0] PE_wrapper207_U0_fifo_w_out_V_V_din_pass_0_out;
  wire fifo_w_PE_4_10_V_V_full_n_pass_0_in;
  wire PE_wrapper207_U0_fifo_w_out_V_V_write_pass_0_out;
  wire [31:0] PE_wrapper183_U0_fifo_cout_drain_out_V_din_pass_0_in;
  wire fifo_cout_drain_PE_2_9_V_full_n_pass_0_out;
  wire PE_wrapper183_U0_fifo_cout_drain_out_V_write_pass_0_in;
  wire [63:0] cout_drain_IO_L1_out_wrapper522_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_9_4_V_V_full_n_pass_0_in;
  wire cout_drain_IO_L1_out_wrapper522_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  wire [63:0] cout_drain_IO_L1_out_wrapper540_U0_fifo_cout_drain_out_V_V_din_pass_0_in;
  wire fifo_cout_drain_cout_drain_IO_L1_out_10_2_V_V_full_n_pass_0_out;
  wire cout_drain_IO_L1_out_wrapper540_U0_fifo_cout_drain_out_V_V_write_pass_0_in;
  wire [63:0] cout_drain_IO_L1_out_wrapper542_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_10_0_V_V_full_n_pass_0_in;
  wire cout_drain_IO_L1_out_wrapper542_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper219_U0_fifo_cin_out_V_V_din_pass_0_out;
  wire fifo_cin_PE_6_9_V_V_full_n_pass_0_in;
  wire PE_wrapper219_U0_fifo_cin_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper172_U0_fifo_cin_out_V_V_din_pass_0_out;
  wire fifo_cin_PE_2_10_V_V_full_n_pass_0_in;
  wire PE_wrapper172_U0_fifo_cin_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper195_U0_fifo_cin_out_V_V_din_pass_1_in;
  wire fifo_cin_PE_4_9_V_V_full_n_pass_1_out;
  wire PE_wrapper195_U0_fifo_cin_out_V_V_write_pass_1_in;
  wire [255:0] cin_IO_L2_in134_U0_fifo_cin_out_V_V_din_pass_0_out;
  wire fifo_cin_cin_IO_L2_in_11_V_V_full_n_pass_0_in;
  wire cin_IO_L2_in134_U0_fifo_cin_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper218_U0_fifo_w_out_V_V_din_pass_0_in;
  wire fifo_w_PE_5_9_V_V_full_n_pass_0_out;
  wire PE_wrapper218_U0_fifo_w_out_V_V_write_pass_0_in;
  wire [63:0] cout_drain_IO_L1_out_wrapper521_U0_fifo_cout_drain_out_V_V_din_pass_1_in;
  wire fifo_cout_drain_cout_drain_IO_L1_out_9_5_V_V_full_n_pass_1_out;
  wire cout_drain_IO_L1_out_wrapper521_U0_fifo_cout_drain_out_V_V_write_pass_1_in;
  wire [31:0] PE_wrapper219_U0_fifo_cout_drain_out_V_din_pass_0_out;
  wire fifo_cout_drain_PE_5_9_V_full_n_pass_0_in;
  wire PE_wrapper219_U0_fifo_cout_drain_out_V_write_pass_0_out;
  wire ap_start_Boundary_X6Y12_To_X8Y12_in;
  wire ap_rst_n_Boundary_X6Y12_To_X8Y12_in;
  wire ap_done_Boundary_X6Y12_To_X8Y12_out;
  wire ap_start_Boundary_X6Y14_To_X8Y14_out;
  wire ap_rst_n_Boundary_X6Y14_To_X8Y14_out;
  wire ap_done_Boundary_X6Y14_To_X8Y14_in;
  wire [255:0] PE_wrapper231_U0_fifo_cin_out_V_V_din_pass_0_in;
  wire [255:0] PE_wrapper231_U0_fifo_cin_out_V_V_din_pass_1_out;
  wire fifo_cin_PE_7_9_V_V_full_n_pass_0_out;
  wire fifo_cin_PE_7_9_V_V_full_n_pass_1_in;
  wire PE_wrapper231_U0_fifo_cin_out_V_V_write_pass_0_in;
  wire PE_wrapper231_U0_fifo_cin_out_V_V_write_pass_1_out;
  wire [63:0] cout_drain_IO_L1_out_wrapper523_U0_fifo_cout_drain_out_V_V_din_pass_0_in;
  wire [63:0] cout_drain_IO_L1_out_wrapper523_U0_fifo_cout_drain_out_V_V_din_pass_1_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_9_3_V_V_full_n_pass_0_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_9_3_V_V_full_n_pass_1_in;
  wire cout_drain_IO_L1_out_wrapper523_U0_fifo_cout_drain_out_V_V_write_pass_0_in;
  wire cout_drain_IO_L1_out_wrapper523_U0_fifo_cout_drain_out_V_V_write_pass_1_out;
  wire [63:0] cout_drain_IO_L2_out558_U0_fifo_cout_drain_out_V_V_din_pass_0_in;
  wire [63:0] cout_drain_IO_L2_out558_U0_fifo_cout_drain_out_V_V_din_pass_1_out;
  wire fifo_cout_drain_cout_drain_IO_L2_out_10_V_V_full_n_pass_0_out;
  wire fifo_cout_drain_cout_drain_IO_L2_out_10_V_V_full_n_pass_1_in;
  wire cout_drain_IO_L2_out558_U0_fifo_cout_drain_out_V_V_write_pass_0_in;
  wire cout_drain_IO_L2_out558_U0_fifo_cout_drain_out_V_V_write_pass_1_out;
  wire [255:0] PE_wrapper195_U0_fifo_cin_out_V_V_din_pass_0_in;
  wire [255:0] PE_wrapper195_U0_fifo_cin_out_V_V_din_pass_1_out;
  wire fifo_cin_PE_4_9_V_V_full_n_pass_0_out;
  wire fifo_cin_PE_4_9_V_V_full_n_pass_1_in;
  wire PE_wrapper195_U0_fifo_cin_out_V_V_write_pass_0_in;
  wire PE_wrapper195_U0_fifo_cin_out_V_V_write_pass_1_out;
  wire [63:0] cout_drain_IO_L1_out_wrapper521_U0_fifo_cout_drain_out_V_V_din_pass_0_in;
  wire [63:0] cout_drain_IO_L1_out_wrapper521_U0_fifo_cout_drain_out_V_V_din_pass_1_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_9_5_V_V_full_n_pass_0_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_9_5_V_V_full_n_pass_1_in;
  wire cout_drain_IO_L1_out_wrapper521_U0_fifo_cout_drain_out_V_V_write_pass_0_in;
  wire cout_drain_IO_L1_out_wrapper521_U0_fifo_cout_drain_out_V_V_write_pass_1_out;
  wire [63:0] cout_drain_IO_L1_out_wrapper551_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_11_6_V_V_full_n_pass_0_in;
  wire cout_drain_IO_L1_out_wrapper551_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  wire [63:0] cout_drain_IO_L1_out_wrapper556_U0_fifo_cout_drain_out_V_V_din_pass_0_in;
  wire fifo_cout_drain_cout_drain_IO_L1_out_11_1_V_V_full_n_pass_0_out;
  wire cout_drain_IO_L1_out_wrapper556_U0_fifo_cout_drain_out_V_V_write_pass_0_in;
  wire [255:0] PE_wrapper160_U0_fifo_w_out_V_V_din_pass_0_in;
  wire fifo_w_PE_0_11_V_V_full_n_pass_0_out;
  wire PE_wrapper160_U0_fifo_w_out_V_V_write_pass_0_in;
  wire [255:0] PE_wrapper244_U0_fifo_cin_out_V_V_din_pass_1_in;
  wire fifo_cin_PE_8_10_V_V_full_n_pass_1_out;
  wire PE_wrapper244_U0_fifo_cin_out_V_V_write_pass_1_in;
  wire [255:0] PE_wrapper173_U0_fifo_w_out_V_V_din_pass_1_in;
  wire fifo_w_PE_1_12_V_V_full_n_pass_1_out;
  wire PE_wrapper173_U0_fifo_w_out_V_V_write_pass_1_in;
  wire [255:0] PE_wrapper184_U0_fifo_w_out_V_V_din_pass_0_in;
  wire fifo_w_PE_2_11_V_V_full_n_pass_0_out;
  wire PE_wrapper184_U0_fifo_w_out_V_V_write_pass_0_in;
  wire [255:0] PE_wrapper161_U0_fifo_cin_out_V_V_din_pass_0_out;
  wire fifo_cin_PE_1_11_V_V_full_n_pass_0_in;
  wire PE_wrapper161_U0_fifo_cin_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper256_U0_fifo_cin_out_V_V_din_pass_0_out;
  wire fifo_cin_PE_9_10_V_V_full_n_pass_0_in;
  wire PE_wrapper256_U0_fifo_cin_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper196_U0_fifo_w_out_V_V_din_pass_0_in;
  wire fifo_w_PE_3_11_V_V_full_n_pass_0_out;
  wire PE_wrapper196_U0_fifo_w_out_V_V_write_pass_0_in;
  wire [255:0] PE_wrapper209_U0_fifo_w_out_V_V_din_pass_0_in;
  wire fifo_w_PE_4_12_V_V_full_n_pass_0_out;
  wire PE_wrapper209_U0_fifo_w_out_V_V_write_pass_0_in;
  wire [255:0] PE_wrapper233_U0_fifo_cin_out_V_V_din_pass_0_in;
  wire fifo_cin_PE_7_11_V_V_full_n_pass_0_out;
  wire PE_wrapper233_U0_fifo_cin_out_V_V_write_pass_0_in;
  wire [31:0] PE_wrapper255_U0_fifo_cout_drain_out_V_din_pass_1_in;
  wire fifo_cout_drain_PE_8_9_V_full_n_pass_1_out;
  wire PE_wrapper255_U0_fifo_cout_drain_out_V_write_pass_1_in;
  wire [255:0] PE_wrapper197_U0_fifo_cin_out_V_V_din_pass_0_out;
  wire fifo_cin_PE_4_11_V_V_full_n_pass_0_in;
  wire PE_wrapper197_U0_fifo_cin_out_V_V_write_pass_0_out;
  wire [31:0] PE_wrapper185_U0_fifo_cout_drain_out_V_din_pass_0_out;
  wire fifo_cout_drain_PE_2_11_V_full_n_pass_0_in;
  wire PE_wrapper185_U0_fifo_cout_drain_out_V_write_pass_0_out;
  wire [63:0] cout_drain_IO_L1_out_wrapper518_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_9_8_V_V_full_n_pass_0_in;
  wire cout_drain_IO_L1_out_wrapper518_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper244_U0_fifo_w_out_V_V_din_pass_1_in;
  wire fifo_w_PE_7_11_V_V_full_n_pass_1_out;
  wire PE_wrapper244_U0_fifo_w_out_V_V_write_pass_1_in;
  wire [63:0] cout_drain_IO_L1_out_wrapper517_U0_fifo_cout_drain_out_V_V_din_pass_2_in;
  wire fifo_cout_drain_cout_drain_IO_L1_out_9_9_V_V_full_n_pass_2_out;
  wire cout_drain_IO_L1_out_wrapper517_U0_fifo_cout_drain_out_V_V_write_pass_2_in;
  wire [63:0] cout_drain_IO_L1_out_wrapper549_U0_fifo_cout_drain_out_V_V_din_pass_0_in;
  wire fifo_cout_drain_cout_drain_IO_L1_out_11_8_V_V_full_n_pass_0_out;
  wire cout_drain_IO_L1_out_wrapper549_U0_fifo_cout_drain_out_V_V_write_pass_0_in;
  wire [255:0] PE_wrapper255_U0_fifo_w_out_V_V_din_pass_1_in;
  wire fifo_w_PE_8_10_V_V_full_n_pass_1_out;
  wire PE_wrapper255_U0_fifo_w_out_V_V_write_pass_1_in;
  wire [63:0] cout_drain_IO_L1_out_wrapper534_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  wire fifo_cout_drain_cout_drain_IO_L1_out_10_8_V_V_full_n_pass_0_in;
  wire cout_drain_IO_L1_out_wrapper534_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  wire [255:0] PE_wrapper257_U0_fifo_cin_out_V_V_din_pass_0_out;
  wire fifo_cin_PE_9_11_V_V_full_n_pass_0_in;
  wire PE_wrapper257_U0_fifo_cin_out_V_V_write_pass_0_out;
  wire [31:0] PE_wrapper257_U0_fifo_cout_drain_out_V_din_pass_0_out;
  wire fifo_cout_drain_PE_8_11_V_full_n_pass_0_in;
  wire PE_wrapper257_U0_fifo_cout_drain_out_V_write_pass_0_out;
  wire [255:0] cin_IO_L2_in_boundary_U0_fifo_cin_local_out_V_V_din_pass_0_in;
  wire fifo_cin_PE_0_11_V_V_full_n_pass_0_out;
  wire cin_IO_L2_in_boundary_U0_fifo_cin_local_out_V_V_write_pass_0_in;
  wire [255:0] PE_wrapper173_U0_fifo_cin_out_V_V_din_pass_1_in;
  wire fifo_cin_PE_2_11_V_V_full_n_pass_1_out;
  wire PE_wrapper173_U0_fifo_cin_out_V_V_write_pass_1_in;
  wire [63:0] cout_drain_IO_L1_out_wrapper533_U0_fifo_cout_drain_out_V_V_din_pass_2_in;
  wire fifo_cout_drain_cout_drain_IO_L1_out_10_9_V_V_full_n_pass_2_out;
  wire cout_drain_IO_L1_out_wrapper533_U0_fifo_cout_drain_out_V_V_write_pass_2_in;
  wire [31:0] PE_wrapper197_U0_fifo_cout_drain_out_V_din_pass_0_out;
  wire fifo_cout_drain_PE_3_11_V_full_n_pass_0_in;
  wire PE_wrapper197_U0_fifo_cout_drain_out_V_write_pass_0_out;
  wire [31:0] PE_wrapper233_U0_fifo_cout_drain_out_V_din_pass_0_in;
  wire fifo_cout_drain_PE_6_11_V_full_n_pass_0_out;
  wire PE_wrapper233_U0_fifo_cout_drain_out_V_write_pass_0_in;
  wire [255:0] PE_wrapper185_U0_fifo_w_out_V_V_din_pass_0_out;
  wire fifo_w_PE_2_12_V_V_full_n_pass_0_in;
  wire PE_wrapper185_U0_fifo_w_out_V_V_write_pass_0_out;
  wire [63:0] cout_drain_IO_L2_out_boundary_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  wire fifo_cout_drain_cout_drain_IO_L2_out_11_V_V_full_n_pass_0_in;
  wire cout_drain_IO_L2_out_boundary_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  wire ap_start_Boundary_X6Y14_To_X8Y14_in;
  wire ap_rst_n_Boundary_X6Y14_To_X8Y14_in;
  wire ap_done_Boundary_X6Y14_To_X8Y14_out;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper211_U0_fifo_cin_out_V_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper211_U0_fifo_cin_out_V_V_din_pass_1_q0 <= PE_wrapper211_U0_fifo_cin_out_V_V_din_pass_1_out;
  end
  assign PE_wrapper211_U0_fifo_cin_out_V_V_din_pass_1_in = PE_wrapper211_U0_fifo_cin_out_V_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_6_1_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_6_1_V_V_full_n_pass_0_q0 <= fifo_cin_PE_6_1_V_V_full_n_pass_0_out;
  end
  assign fifo_cin_PE_6_1_V_V_full_n_pass_0_in = fifo_cin_PE_6_1_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper211_U0_fifo_cin_out_V_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper211_U0_fifo_cin_out_V_V_write_pass_1_q0 <= PE_wrapper211_U0_fifo_cin_out_V_V_write_pass_1_out;
  end
  assign PE_wrapper211_U0_fifo_cin_out_V_V_write_pass_1_in = PE_wrapper211_U0_fifo_cin_out_V_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper212_U0_fifo_cin_out_V_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper212_U0_fifo_cin_out_V_V_din_pass_1_q0 <= PE_wrapper212_U0_fifo_cin_out_V_V_din_pass_1_out;
  end
  assign PE_wrapper212_U0_fifo_cin_out_V_V_din_pass_1_in = PE_wrapper212_U0_fifo_cin_out_V_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_6_2_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_6_2_V_V_full_n_pass_0_q0 <= fifo_cin_PE_6_2_V_V_full_n_pass_0_out;
  end
  assign fifo_cin_PE_6_2_V_V_full_n_pass_0_in = fifo_cin_PE_6_2_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper212_U0_fifo_cin_out_V_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper212_U0_fifo_cin_out_V_V_write_pass_1_q0 <= PE_wrapper212_U0_fifo_cin_out_V_V_write_pass_1_out;
  end
  assign PE_wrapper212_U0_fifo_cin_out_V_V_write_pass_1_in = PE_wrapper212_U0_fifo_cin_out_V_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper213_U0_fifo_cin_out_V_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper213_U0_fifo_cin_out_V_V_din_pass_1_q0 <= PE_wrapper213_U0_fifo_cin_out_V_V_din_pass_1_out;
  end
  assign PE_wrapper213_U0_fifo_cin_out_V_V_din_pass_1_in = PE_wrapper213_U0_fifo_cin_out_V_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_6_3_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_6_3_V_V_full_n_pass_0_q0 <= fifo_cin_PE_6_3_V_V_full_n_pass_0_out;
  end
  assign fifo_cin_PE_6_3_V_V_full_n_pass_0_in = fifo_cin_PE_6_3_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper213_U0_fifo_cin_out_V_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper213_U0_fifo_cin_out_V_V_write_pass_1_q0 <= PE_wrapper213_U0_fifo_cin_out_V_V_write_pass_1_out;
  end
  assign PE_wrapper213_U0_fifo_cin_out_V_V_write_pass_1_in = PE_wrapper213_U0_fifo_cin_out_V_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [255:0] cin_IO_L2_in125_U0_fifo_cin_out_V_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    cin_IO_L2_in125_U0_fifo_cin_out_V_V_din_pass_1_q0 <= cin_IO_L2_in125_U0_fifo_cin_out_V_V_din_pass_1_out;
  end
  assign cin_IO_L2_in125_U0_fifo_cin_out_V_V_din_pass_1_in = cin_IO_L2_in125_U0_fifo_cin_out_V_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_cin_IO_L2_in_2_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_cin_IO_L2_in_2_V_V_full_n_pass_0_q0 <= fifo_cin_cin_IO_L2_in_2_V_V_full_n_pass_0_out;
  end
  assign fifo_cin_cin_IO_L2_in_2_V_V_full_n_pass_0_in = fifo_cin_cin_IO_L2_in_2_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  cin_IO_L2_in125_U0_fifo_cin_out_V_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    cin_IO_L2_in125_U0_fifo_cin_out_V_V_write_pass_1_q0 <= cin_IO_L2_in125_U0_fifo_cin_out_V_V_write_pass_1_out;
  end
  assign cin_IO_L2_in125_U0_fifo_cin_out_V_V_write_pass_1_in = cin_IO_L2_in125_U0_fifo_cin_out_V_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [63:0] cout_drain_IO_L1_out_wrapper424_U0_fifo_cout_drain_out_V_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper424_U0_fifo_cout_drain_out_V_V_din_pass_1_q0 <= cout_drain_IO_L1_out_wrapper424_U0_fifo_cout_drain_out_V_V_din_pass_1_out;
  end
  assign cout_drain_IO_L1_out_wrapper424_U0_fifo_cout_drain_out_V_V_din_pass_1_in = cout_drain_IO_L1_out_wrapper424_U0_fifo_cout_drain_out_V_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_cout_drain_IO_L1_out_3_6_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_cout_drain_IO_L1_out_3_6_V_V_full_n_pass_0_q0 <= fifo_cout_drain_cout_drain_IO_L1_out_3_6_V_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_cout_drain_IO_L1_out_3_6_V_V_full_n_pass_0_in = fifo_cout_drain_cout_drain_IO_L1_out_3_6_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  cout_drain_IO_L1_out_wrapper424_U0_fifo_cout_drain_out_V_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper424_U0_fifo_cout_drain_out_V_V_write_pass_1_q0 <= cout_drain_IO_L1_out_wrapper424_U0_fifo_cout_drain_out_V_V_write_pass_1_out;
  end
  assign cout_drain_IO_L1_out_wrapper424_U0_fifo_cout_drain_out_V_V_write_pass_1_in = cout_drain_IO_L1_out_wrapper424_U0_fifo_cout_drain_out_V_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [63:0] cout_drain_IO_L1_out_wrapper408_U0_fifo_cout_drain_out_V_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper408_U0_fifo_cout_drain_out_V_V_din_pass_1_q0 <= cout_drain_IO_L1_out_wrapper408_U0_fifo_cout_drain_out_V_V_din_pass_1_out;
  end
  assign cout_drain_IO_L1_out_wrapper408_U0_fifo_cout_drain_out_V_V_din_pass_1_in = cout_drain_IO_L1_out_wrapper408_U0_fifo_cout_drain_out_V_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_cout_drain_IO_L1_out_2_6_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_cout_drain_IO_L1_out_2_6_V_V_full_n_pass_0_q0 <= fifo_cout_drain_cout_drain_IO_L1_out_2_6_V_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_cout_drain_IO_L1_out_2_6_V_V_full_n_pass_0_in = fifo_cout_drain_cout_drain_IO_L1_out_2_6_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  cout_drain_IO_L1_out_wrapper408_U0_fifo_cout_drain_out_V_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper408_U0_fifo_cout_drain_out_V_V_write_pass_1_q0 <= cout_drain_IO_L1_out_wrapper408_U0_fifo_cout_drain_out_V_V_write_pass_1_out;
  end
  assign cout_drain_IO_L1_out_wrapper408_U0_fifo_cout_drain_out_V_V_write_pass_1_in = cout_drain_IO_L1_out_wrapper408_U0_fifo_cout_drain_out_V_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [63:0] cout_drain_IO_L1_out_wrapper376_U0_fifo_cout_drain_out_V_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper376_U0_fifo_cout_drain_out_V_V_din_pass_1_q0 <= cout_drain_IO_L1_out_wrapper376_U0_fifo_cout_drain_out_V_V_din_pass_1_out;
  end
  assign cout_drain_IO_L1_out_wrapper376_U0_fifo_cout_drain_out_V_V_din_pass_1_in = cout_drain_IO_L1_out_wrapper376_U0_fifo_cout_drain_out_V_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_cout_drain_IO_L1_out_0_6_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_cout_drain_IO_L1_out_0_6_V_V_full_n_pass_0_q0 <= fifo_cout_drain_cout_drain_IO_L1_out_0_6_V_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_cout_drain_IO_L1_out_0_6_V_V_full_n_pass_0_in = fifo_cout_drain_cout_drain_IO_L1_out_0_6_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  cout_drain_IO_L1_out_wrapper376_U0_fifo_cout_drain_out_V_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper376_U0_fifo_cout_drain_out_V_V_write_pass_1_q0 <= cout_drain_IO_L1_out_wrapper376_U0_fifo_cout_drain_out_V_V_write_pass_1_out;
  end
  assign cout_drain_IO_L1_out_wrapper376_U0_fifo_cout_drain_out_V_V_write_pass_1_in = cout_drain_IO_L1_out_wrapper376_U0_fifo_cout_drain_out_V_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [63:0] cout_drain_IO_L1_out_wrapper392_U0_fifo_cout_drain_out_V_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper392_U0_fifo_cout_drain_out_V_V_din_pass_1_q0 <= cout_drain_IO_L1_out_wrapper392_U0_fifo_cout_drain_out_V_V_din_pass_1_out;
  end
  assign cout_drain_IO_L1_out_wrapper392_U0_fifo_cout_drain_out_V_V_din_pass_1_in = cout_drain_IO_L1_out_wrapper392_U0_fifo_cout_drain_out_V_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_cout_drain_IO_L1_out_1_6_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_cout_drain_IO_L1_out_1_6_V_V_full_n_pass_0_q0 <= fifo_cout_drain_cout_drain_IO_L1_out_1_6_V_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_cout_drain_IO_L1_out_1_6_V_V_full_n_pass_0_in = fifo_cout_drain_cout_drain_IO_L1_out_1_6_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  cout_drain_IO_L1_out_wrapper392_U0_fifo_cout_drain_out_V_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper392_U0_fifo_cout_drain_out_V_V_write_pass_1_q0 <= cout_drain_IO_L1_out_wrapper392_U0_fifo_cout_drain_out_V_V_write_pass_1_out;
  end
  assign cout_drain_IO_L1_out_wrapper392_U0_fifo_cout_drain_out_V_V_write_pass_1_in = cout_drain_IO_L1_out_wrapper392_U0_fifo_cout_drain_out_V_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper213_U0_fifo_w_out_V_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper213_U0_fifo_w_out_V_V_din_pass_1_q0 <= PE_wrapper213_U0_fifo_w_out_V_V_din_pass_1_out;
  end
  assign PE_wrapper213_U0_fifo_w_out_V_V_din_pass_1_in = PE_wrapper213_U0_fifo_w_out_V_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_5_4_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_5_4_V_V_full_n_pass_0_q0 <= fifo_w_PE_5_4_V_V_full_n_pass_0_out;
  end
  assign fifo_w_PE_5_4_V_V_full_n_pass_0_in = fifo_w_PE_5_4_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper213_U0_fifo_w_out_V_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper213_U0_fifo_w_out_V_V_write_pass_1_q0 <= PE_wrapper213_U0_fifo_w_out_V_V_write_pass_1_out;
  end
  assign PE_wrapper213_U0_fifo_w_out_V_V_write_pass_1_in = PE_wrapper213_U0_fifo_w_out_V_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper187_U0_fifo_w_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper187_U0_fifo_w_out_V_V_din_pass_0_q0 <= PE_wrapper187_U0_fifo_w_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper187_U0_fifo_w_out_V_V_din_pass_0_in = PE_wrapper187_U0_fifo_w_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper187_U0_fifo_w_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper187_U0_fifo_w_out_V_V_write_pass_0_q0 <= PE_wrapper187_U0_fifo_w_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper187_U0_fifo_w_out_V_V_write_pass_0_in = PE_wrapper187_U0_fifo_w_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [31:0] PE_wrapper187_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper187_U0_fifo_cout_drain_out_V_din_pass_0_q0 <= PE_wrapper187_U0_fifo_cout_drain_out_V_din_pass_0_out;
  end
  assign PE_wrapper187_U0_fifo_cout_drain_out_V_din_pass_0_in = PE_wrapper187_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper187_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper187_U0_fifo_cout_drain_out_V_write_pass_0_q0 <= PE_wrapper187_U0_fifo_cout_drain_out_V_write_pass_0_out;
  end
  assign PE_wrapper187_U0_fifo_cout_drain_out_V_write_pass_0_in = PE_wrapper187_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_2_0_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_2_0_V_V_full_n_pass_0_q0 <= fifo_cin_PE_2_0_V_V_full_n_pass_0_out;
  end
  assign fifo_cin_PE_2_0_V_V_full_n_pass_0_in = fifo_cin_PE_2_0_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] w_IO_L2_in137_U0_fifo_w_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    w_IO_L2_in137_U0_fifo_w_out_V_V_din_pass_0_q0 <= w_IO_L2_in137_U0_fifo_w_out_V_V_din_pass_0_out;
  end
  assign w_IO_L2_in137_U0_fifo_w_out_V_V_din_pass_0_in = w_IO_L2_in137_U0_fifo_w_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  w_IO_L2_in137_U0_fifo_w_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    w_IO_L2_in137_U0_fifo_w_out_V_V_write_pass_0_q0 <= w_IO_L2_in137_U0_fifo_w_out_V_V_write_pass_0_out;
  end
  assign w_IO_L2_in137_U0_fifo_w_out_V_V_write_pass_0_in = w_IO_L2_in137_U0_fifo_w_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [31:0] PE_wrapper151_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper151_U0_fifo_cout_drain_out_V_din_pass_0_q0 <= PE_wrapper151_U0_fifo_cout_drain_out_V_din_pass_0_out;
  end
  assign PE_wrapper151_U0_fifo_cout_drain_out_V_din_pass_0_in = PE_wrapper151_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper151_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper151_U0_fifo_cout_drain_out_V_write_pass_0_q0 <= PE_wrapper151_U0_fifo_cout_drain_out_V_write_pass_0_out;
  end
  assign PE_wrapper151_U0_fifo_cout_drain_out_V_write_pass_0_in = PE_wrapper151_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper163_U0_fifo_w_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper163_U0_fifo_w_out_V_V_din_pass_0_q0 <= PE_wrapper163_U0_fifo_w_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper163_U0_fifo_w_out_V_V_din_pass_0_in = PE_wrapper163_U0_fifo_w_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper163_U0_fifo_w_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper163_U0_fifo_w_out_V_V_write_pass_0_q0 <= PE_wrapper163_U0_fifo_w_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper163_U0_fifo_w_out_V_V_write_pass_0_in = PE_wrapper163_U0_fifo_w_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_w_w_IO_L2_in_2_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_w_IO_L2_in_2_V_V_full_n_pass_0_q0 <= fifo_w_w_IO_L2_in_2_V_V_full_n_pass_0_out;
  end
  assign fifo_w_w_IO_L2_in_2_V_V_full_n_pass_0_in = fifo_w_w_IO_L2_in_2_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] cin_IO_L2_in124_U0_fifo_cin_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    cin_IO_L2_in124_U0_fifo_cin_out_V_V_din_pass_0_q0 <= cin_IO_L2_in124_U0_fifo_cin_out_V_V_din_pass_0_out;
  end
  assign cin_IO_L2_in124_U0_fifo_cin_out_V_V_din_pass_0_in = cin_IO_L2_in124_U0_fifo_cin_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  cin_IO_L2_in124_U0_fifo_cin_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    cin_IO_L2_in124_U0_fifo_cin_out_V_V_write_pass_0_q0 <= cin_IO_L2_in124_U0_fifo_cin_out_V_V_write_pass_0_out;
  end
  assign cin_IO_L2_in124_U0_fifo_cin_out_V_V_write_pass_0_in = cin_IO_L2_in124_U0_fifo_cin_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_3_0_V_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_3_0_V_V_full_n_pass_1_q0 <= fifo_w_PE_3_0_V_V_full_n_pass_1_out;
  end
  assign fifo_w_PE_3_0_V_V_full_n_pass_1_in = fifo_w_PE_3_0_V_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg [63:0] kernel0_entry12_U0_w_V_out_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    kernel0_entry12_U0_w_V_out_din_pass_0_q0 <= kernel0_entry12_U0_w_V_out_din_pass_0_out;
  end
  assign kernel0_entry12_U0_w_V_out_din_pass_0_in = kernel0_entry12_U0_w_V_out_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  kernel0_entry12_U0_w_V_out_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    kernel0_entry12_U0_w_V_out_write_pass_0_q0 <= kernel0_entry12_U0_w_V_out_write_pass_0_out;
  end
  assign kernel0_entry12_U0_w_V_out_write_pass_0_in = kernel0_entry12_U0_w_V_out_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [31:0] PE_wrapper163_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper163_U0_fifo_cout_drain_out_V_din_pass_0_q0 <= PE_wrapper163_U0_fifo_cout_drain_out_V_din_pass_0_out;
  end
  assign PE_wrapper163_U0_fifo_cout_drain_out_V_din_pass_0_in = PE_wrapper163_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper163_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper163_U0_fifo_cout_drain_out_V_write_pass_0_q0 <= PE_wrapper163_U0_fifo_cout_drain_out_V_write_pass_0_out;
  end
  assign PE_wrapper163_U0_fifo_cout_drain_out_V_write_pass_0_in = PE_wrapper163_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper151_U0_fifo_w_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper151_U0_fifo_w_out_V_V_din_pass_0_q0 <= PE_wrapper151_U0_fifo_w_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper151_U0_fifo_w_out_V_V_din_pass_0_in = PE_wrapper151_U0_fifo_w_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper151_U0_fifo_w_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper151_U0_fifo_w_out_V_V_write_pass_0_q0 <= PE_wrapper151_U0_fifo_w_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper151_U0_fifo_w_out_V_V_write_pass_0_in = PE_wrapper151_U0_fifo_w_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_PE_1_0_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_PE_1_0_V_full_n_pass_0_q0 <= fifo_cout_drain_PE_1_0_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_PE_1_0_V_full_n_pass_0_in = fifo_cout_drain_PE_1_0_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper150_U0_fifo_cin_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper150_U0_fifo_cin_out_V_V_din_pass_0_q0 <= PE_wrapper150_U0_fifo_cin_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper150_U0_fifo_cin_out_V_V_din_pass_0_in = PE_wrapper150_U0_fifo_cin_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper150_U0_fifo_cin_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper150_U0_fifo_cin_out_V_V_write_pass_0_q0 <= PE_wrapper150_U0_fifo_cin_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper150_U0_fifo_cin_out_V_V_write_pass_0_in = PE_wrapper150_U0_fifo_cin_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [31:0] PE_wrapper175_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper175_U0_fifo_cout_drain_out_V_din_pass_0_q0 <= PE_wrapper175_U0_fifo_cout_drain_out_V_din_pass_0_out;
  end
  assign PE_wrapper175_U0_fifo_cout_drain_out_V_din_pass_0_in = PE_wrapper175_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper175_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper175_U0_fifo_cout_drain_out_V_write_pass_0_q0 <= PE_wrapper175_U0_fifo_cout_drain_out_V_write_pass_0_out;
  end
  assign PE_wrapper175_U0_fifo_cout_drain_out_V_write_pass_0_in = PE_wrapper175_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper175_U0_fifo_w_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper175_U0_fifo_w_out_V_V_din_pass_0_q0 <= PE_wrapper175_U0_fifo_w_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper175_U0_fifo_w_out_V_V_din_pass_0_in = PE_wrapper175_U0_fifo_w_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper175_U0_fifo_w_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper175_U0_fifo_w_out_V_V_write_pass_0_q0 <= PE_wrapper175_U0_fifo_w_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper175_U0_fifo_w_out_V_V_write_pass_0_in = PE_wrapper175_U0_fifo_w_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_0_1_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_0_1_V_V_full_n_pass_0_q0 <= fifo_cin_PE_0_1_V_V_full_n_pass_0_out;
  end
  assign fifo_cin_PE_0_1_V_V_full_n_pass_0_in = fifo_cin_PE_0_1_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_cout_drain_IO_L1_out_0_4_V_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_cout_drain_IO_L1_out_0_4_V_V_full_n_pass_1_q0 <= fifo_cout_drain_cout_drain_IO_L1_out_0_4_V_V_full_n_pass_1_out;
  end
  assign fifo_cout_drain_cout_drain_IO_L1_out_0_4_V_V_full_n_pass_1_in = fifo_cout_drain_cout_drain_IO_L1_out_0_4_V_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg [63:0] kernel0_entry12_U0_cout_V_out_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    kernel0_entry12_U0_cout_V_out_din_pass_0_q0 <= kernel0_entry12_U0_cout_V_out_din_pass_0_out;
  end
  assign kernel0_entry12_U0_cout_V_out_din_pass_0_in = kernel0_entry12_U0_cout_V_out_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  kernel0_entry12_U0_cout_V_out_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    kernel0_entry12_U0_cout_V_out_write_pass_0_q0 <= kernel0_entry12_U0_cout_V_out_write_pass_0_out;
  end
  assign kernel0_entry12_U0_cout_V_out_write_pass_0_in = kernel0_entry12_U0_cout_V_out_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper187_U0_fifo_cin_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper187_U0_fifo_cin_out_V_V_din_pass_0_q0 <= PE_wrapper187_U0_fifo_cin_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper187_U0_fifo_cin_out_V_V_din_pass_0_in = PE_wrapper187_U0_fifo_cin_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper187_U0_fifo_cin_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper187_U0_fifo_cin_out_V_V_write_pass_0_q0 <= PE_wrapper187_U0_fifo_cin_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper187_U0_fifo_cin_out_V_V_write_pass_0_in = PE_wrapper187_U0_fifo_cin_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_1_1_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_1_1_V_V_full_n_pass_0_q0 <= fifo_w_PE_1_1_V_V_full_n_pass_0_out;
  end
  assign fifo_w_PE_1_1_V_V_full_n_pass_0_in = fifo_w_PE_1_1_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg [63:0] cout_drain_IO_L1_out_wrapper382_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper382_U0_fifo_cout_drain_out_V_V_din_pass_0_q0 <= cout_drain_IO_L1_out_wrapper382_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper382_U0_fifo_cout_drain_out_V_V_din_pass_0_in = cout_drain_IO_L1_out_wrapper382_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  cout_drain_IO_L1_out_wrapper382_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper382_U0_fifo_cout_drain_out_V_V_write_pass_0_q0 <= cout_drain_IO_L1_out_wrapper382_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper382_U0_fifo_cout_drain_out_V_V_write_pass_0_in = cout_drain_IO_L1_out_wrapper382_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper186_U0_fifo_cin_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper186_U0_fifo_cin_out_V_V_din_pass_0_q0 <= PE_wrapper186_U0_fifo_cin_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper186_U0_fifo_cin_out_V_V_din_pass_0_in = PE_wrapper186_U0_fifo_cin_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper186_U0_fifo_cin_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper186_U0_fifo_cin_out_V_V_write_pass_0_q0 <= PE_wrapper186_U0_fifo_cin_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper186_U0_fifo_cin_out_V_V_write_pass_0_in = PE_wrapper186_U0_fifo_cin_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_0_0_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_0_0_V_V_full_n_pass_0_q0 <= fifo_w_PE_0_0_V_V_full_n_pass_0_out;
  end
  assign fifo_w_PE_0_0_V_V_full_n_pass_0_in = fifo_w_PE_0_0_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  ap_start_Boundary_X4Y2_To_X6Y2_q0;
  always @ (posedge ap_clk) begin
    ap_start_Boundary_X4Y2_To_X6Y2_q0 <= ap_start_Boundary_X4Y2_To_X6Y2_out;
  end
  assign ap_start_Boundary_X4Y2_To_X6Y2_in = ap_start_Boundary_X4Y2_To_X6Y2_q0;
  (* dont_touch = "yes" *) reg  ap_rst_n_Boundary_X4Y2_To_X6Y2_q0;
  always @ (posedge ap_clk) begin
    ap_rst_n_Boundary_X4Y2_To_X6Y2_q0 <= ap_rst_n_Boundary_X4Y2_To_X6Y2_out;
  end
  assign ap_rst_n_Boundary_X4Y2_To_X6Y2_in = ap_rst_n_Boundary_X4Y2_To_X6Y2_q0;
  (* dont_touch = "yes" *) reg  ap_start_Boundary_X6Y0_To_X6Y2_q0;
  always @ (posedge ap_clk) begin
    ap_start_Boundary_X6Y0_To_X6Y2_q0 <= ap_start_Boundary_X6Y0_To_X6Y2_out;
  end
  assign ap_start_Boundary_X6Y0_To_X6Y2_in = ap_start_Boundary_X6Y0_To_X6Y2_q0;
  (* dont_touch = "yes" *) reg  ap_rst_n_Boundary_X6Y0_To_X6Y2_q0;
  always @ (posedge ap_clk) begin
    ap_rst_n_Boundary_X6Y0_To_X6Y2_q0 <= ap_rst_n_Boundary_X6Y0_To_X6Y2_out;
  end
  assign ap_rst_n_Boundary_X6Y0_To_X6Y2_in = ap_rst_n_Boundary_X6Y0_To_X6Y2_q0;
  (* dont_touch = "yes" *) reg  ap_start_Boundary_X4Y0_To_X4Y2_q0;
  always @ (posedge ap_clk) begin
    ap_start_Boundary_X4Y0_To_X4Y2_q0 <= ap_start_Boundary_X4Y0_To_X4Y2_out;
  end
  assign ap_start_Boundary_X4Y0_To_X4Y2_in = ap_start_Boundary_X4Y0_To_X4Y2_q0;
  (* dont_touch = "yes" *) reg  ap_rst_n_Boundary_X4Y0_To_X4Y2_q0;
  always @ (posedge ap_clk) begin
    ap_rst_n_Boundary_X4Y0_To_X4Y2_q0 <= ap_rst_n_Boundary_X4Y0_To_X4Y2_out;
  end
  assign ap_rst_n_Boundary_X4Y0_To_X4Y2_in = ap_rst_n_Boundary_X4Y0_To_X4Y2_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper190_U0_fifo_w_out_V_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper190_U0_fifo_w_out_V_V_din_pass_1_q0 <= PE_wrapper190_U0_fifo_w_out_V_V_din_pass_1_out;
  end
  assign PE_wrapper190_U0_fifo_w_out_V_V_din_pass_1_in = PE_wrapper190_U0_fifo_w_out_V_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_3_5_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_3_5_V_V_full_n_pass_0_q0 <= fifo_w_PE_3_5_V_V_full_n_pass_0_out;
  end
  assign fifo_w_PE_3_5_V_V_full_n_pass_0_in = fifo_w_PE_3_5_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper190_U0_fifo_w_out_V_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper190_U0_fifo_w_out_V_V_write_pass_1_q0 <= PE_wrapper190_U0_fifo_w_out_V_V_write_pass_1_out;
  end
  assign PE_wrapper190_U0_fifo_w_out_V_V_write_pass_1_in = PE_wrapper190_U0_fifo_w_out_V_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper179_U0_fifo_cin_out_V_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper179_U0_fifo_cin_out_V_V_din_pass_1_q0 <= PE_wrapper179_U0_fifo_cin_out_V_V_din_pass_1_out;
  end
  assign PE_wrapper179_U0_fifo_cin_out_V_V_din_pass_1_in = PE_wrapper179_U0_fifo_cin_out_V_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_3_5_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_3_5_V_V_full_n_pass_0_q0 <= fifo_cin_PE_3_5_V_V_full_n_pass_0_out;
  end
  assign fifo_cin_PE_3_5_V_V_full_n_pass_0_in = fifo_cin_PE_3_5_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper179_U0_fifo_cin_out_V_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper179_U0_fifo_cin_out_V_V_write_pass_1_q0 <= PE_wrapper179_U0_fifo_cin_out_V_V_write_pass_1_out;
  end
  assign PE_wrapper179_U0_fifo_cin_out_V_V_write_pass_1_in = PE_wrapper179_U0_fifo_cin_out_V_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [63:0] kernel0_entry12_U0_cout_V_out_din_pass_2_q0;
  always @ (posedge ap_clk) begin
    kernel0_entry12_U0_cout_V_out_din_pass_2_q0 <= kernel0_entry12_U0_cout_V_out_din_pass_2_out;
  end
  assign kernel0_entry12_U0_cout_V_out_din_pass_2_in = kernel0_entry12_U0_cout_V_out_din_pass_2_q0;
  (* dont_touch = "yes" *) reg  cout_V_c_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    cout_V_c_full_n_pass_1_q0 <= cout_V_c_full_n_pass_1_out;
  end
  assign cout_V_c_full_n_pass_1_in = cout_V_c_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg  kernel0_entry12_U0_cout_V_out_write_pass_2_q0;
  always @ (posedge ap_clk) begin
    kernel0_entry12_U0_cout_V_out_write_pass_2_q0 <= kernel0_entry12_U0_cout_V_out_write_pass_2_out;
  end
  assign kernel0_entry12_U0_cout_V_out_write_pass_2_in = kernel0_entry12_U0_cout_V_out_write_pass_2_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_4_4_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_4_4_V_V_full_n_pass_0_q0 <= fifo_cin_PE_4_4_V_V_full_n_pass_0_out;
  end
  assign fifo_cin_PE_4_4_V_V_full_n_pass_0_in = fifo_cin_PE_4_4_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_4_4_V_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_4_4_V_V_full_n_pass_1_q0 <= fifo_w_PE_4_4_V_V_full_n_pass_1_out;
  end
  assign fifo_w_PE_4_4_V_V_full_n_pass_1_in = fifo_w_PE_4_4_V_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_cout_drain_IO_L1_out_4_6_V_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_cout_drain_IO_L1_out_4_6_V_V_full_n_pass_1_q0 <= fifo_cout_drain_cout_drain_IO_L1_out_4_6_V_V_full_n_pass_1_out;
  end
  assign fifo_cout_drain_cout_drain_IO_L1_out_4_6_V_V_full_n_pass_1_in = fifo_cout_drain_cout_drain_IO_L1_out_4_6_V_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_5_4_V_V_full_n_pass_2_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_5_4_V_V_full_n_pass_2_q0 <= fifo_w_PE_5_4_V_V_full_n_pass_2_out;
  end
  assign fifo_w_PE_5_4_V_V_full_n_pass_2_in = fifo_w_PE_5_4_V_V_full_n_pass_2_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper214_U0_fifo_w_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper214_U0_fifo_w_out_V_V_din_pass_0_q0 <= PE_wrapper214_U0_fifo_w_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper214_U0_fifo_w_out_V_V_din_pass_0_in = PE_wrapper214_U0_fifo_w_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper214_U0_fifo_w_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper214_U0_fifo_w_out_V_V_write_pass_0_q0 <= PE_wrapper214_U0_fifo_w_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper214_U0_fifo_w_out_V_V_write_pass_0_in = PE_wrapper214_U0_fifo_w_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [63:0] cout_drain_IO_L1_out_wrapper441_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper441_U0_fifo_cout_drain_out_V_V_din_pass_0_q0 <= cout_drain_IO_L1_out_wrapper441_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper441_U0_fifo_cout_drain_out_V_V_din_pass_0_in = cout_drain_IO_L1_out_wrapper441_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  cout_drain_IO_L1_out_wrapper441_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper441_U0_fifo_cout_drain_out_V_V_write_pass_0_q0 <= cout_drain_IO_L1_out_wrapper441_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper441_U0_fifo_cout_drain_out_V_V_write_pass_0_in = cout_drain_IO_L1_out_wrapper441_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] w_IO_L3_in_serialize_U0_fifo_w_local_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    w_IO_L3_in_serialize_U0_fifo_w_local_out_V_V_din_pass_0_q0 <= w_IO_L3_in_serialize_U0_fifo_w_local_out_V_V_din_pass_0_out;
  end
  assign w_IO_L3_in_serialize_U0_fifo_w_local_out_V_V_din_pass_0_in = w_IO_L3_in_serialize_U0_fifo_w_local_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  w_IO_L3_in_serialize_U0_fifo_w_local_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    w_IO_L3_in_serialize_U0_fifo_w_local_out_V_V_write_pass_0_q0 <= w_IO_L3_in_serialize_U0_fifo_w_local_out_V_V_write_pass_0_out;
  end
  assign w_IO_L3_in_serialize_U0_fifo_w_local_out_V_V_write_pass_0_in = w_IO_L3_in_serialize_U0_fifo_w_local_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper214_U0_fifo_cin_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper214_U0_fifo_cin_out_V_V_din_pass_0_q0 <= PE_wrapper214_U0_fifo_cin_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper214_U0_fifo_cin_out_V_V_din_pass_0_in = PE_wrapper214_U0_fifo_cin_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper214_U0_fifo_cin_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper214_U0_fifo_cin_out_V_V_write_pass_0_q0 <= PE_wrapper214_U0_fifo_cin_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper214_U0_fifo_cin_out_V_V_write_pass_0_in = PE_wrapper214_U0_fifo_cin_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper202_U0_fifo_w_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper202_U0_fifo_w_out_V_V_din_pass_0_q0 <= PE_wrapper202_U0_fifo_w_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper202_U0_fifo_w_out_V_V_din_pass_0_in = PE_wrapper202_U0_fifo_w_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper202_U0_fifo_w_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper202_U0_fifo_w_out_V_V_write_pass_0_q0 <= PE_wrapper202_U0_fifo_w_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper202_U0_fifo_w_out_V_V_write_pass_0_in = PE_wrapper202_U0_fifo_w_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [31:0] PE_wrapper202_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper202_U0_fifo_cout_drain_out_V_din_pass_0_q0 <= PE_wrapper202_U0_fifo_cout_drain_out_V_din_pass_0_out;
  end
  assign PE_wrapper202_U0_fifo_cout_drain_out_V_din_pass_0_in = PE_wrapper202_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper202_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper202_U0_fifo_cout_drain_out_V_write_pass_0_q0 <= PE_wrapper202_U0_fifo_cout_drain_out_V_write_pass_0_out;
  end
  assign PE_wrapper202_U0_fifo_cout_drain_out_V_write_pass_0_in = PE_wrapper202_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  w_V_c_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    w_V_c_full_n_pass_1_q0 <= w_V_c_full_n_pass_1_out;
  end
  assign w_V_c_full_n_pass_1_in = w_V_c_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg  ap_done_Boundary_X4Y4_To_X6Y4_q0;
  always @ (posedge ap_clk) begin
    ap_done_Boundary_X4Y4_To_X6Y4_q0 <= ap_done_Boundary_X4Y4_To_X6Y4_out;
  end
  assign ap_done_Boundary_X4Y4_To_X6Y4_in = ap_done_Boundary_X4Y4_To_X6Y4_q0;
  (* dont_touch = "yes" *) reg  ap_start_Boundary_X4Y6_To_X6Y6_q0;
  always @ (posedge ap_clk) begin
    ap_start_Boundary_X4Y6_To_X6Y6_q0 <= ap_start_Boundary_X4Y6_To_X6Y6_out;
  end
  assign ap_start_Boundary_X4Y6_To_X6Y6_in = ap_start_Boundary_X4Y6_To_X6Y6_q0;
  (* dont_touch = "yes" *) reg  ap_rst_n_Boundary_X4Y6_To_X6Y6_q0;
  always @ (posedge ap_clk) begin
    ap_rst_n_Boundary_X4Y6_To_X6Y6_q0 <= ap_rst_n_Boundary_X4Y6_To_X6Y6_out;
  end
  assign ap_rst_n_Boundary_X4Y6_To_X6Y6_in = ap_rst_n_Boundary_X4Y6_To_X6Y6_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper230_U0_fifo_w_out_V_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper230_U0_fifo_w_out_V_V_din_pass_1_q0 <= PE_wrapper230_U0_fifo_w_out_V_V_din_pass_1_out;
  end
  assign PE_wrapper230_U0_fifo_w_out_V_V_din_pass_1_in = PE_wrapper230_U0_fifo_w_out_V_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_6_9_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_6_9_V_V_full_n_pass_0_q0 <= fifo_w_PE_6_9_V_V_full_n_pass_0_out;
  end
  assign fifo_w_PE_6_9_V_V_full_n_pass_0_in = fifo_w_PE_6_9_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper230_U0_fifo_w_out_V_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper230_U0_fifo_w_out_V_V_write_pass_1_q0 <= PE_wrapper230_U0_fifo_w_out_V_V_write_pass_1_out;
  end
  assign PE_wrapper230_U0_fifo_w_out_V_V_write_pass_1_in = PE_wrapper230_U0_fifo_w_out_V_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [63:0] cout_drain_IO_L1_out_wrapper522_U0_fifo_cout_drain_out_V_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper522_U0_fifo_cout_drain_out_V_V_din_pass_1_q0 <= cout_drain_IO_L1_out_wrapper522_U0_fifo_cout_drain_out_V_V_din_pass_1_out;
  end
  assign cout_drain_IO_L1_out_wrapper522_U0_fifo_cout_drain_out_V_V_din_pass_1_in = cout_drain_IO_L1_out_wrapper522_U0_fifo_cout_drain_out_V_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_cout_drain_IO_L1_out_9_4_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_cout_drain_IO_L1_out_9_4_V_V_full_n_pass_0_q0 <= fifo_cout_drain_cout_drain_IO_L1_out_9_4_V_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_cout_drain_IO_L1_out_9_4_V_V_full_n_pass_0_in = fifo_cout_drain_cout_drain_IO_L1_out_9_4_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  cout_drain_IO_L1_out_wrapper522_U0_fifo_cout_drain_out_V_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper522_U0_fifo_cout_drain_out_V_V_write_pass_1_q0 <= cout_drain_IO_L1_out_wrapper522_U0_fifo_cout_drain_out_V_V_write_pass_1_out;
  end
  assign cout_drain_IO_L1_out_wrapper522_U0_fifo_cout_drain_out_V_V_write_pass_1_in = cout_drain_IO_L1_out_wrapper522_U0_fifo_cout_drain_out_V_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [63:0] cout_drain_IO_L1_out_wrapper542_U0_fifo_cout_drain_out_V_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper542_U0_fifo_cout_drain_out_V_V_din_pass_1_q0 <= cout_drain_IO_L1_out_wrapper542_U0_fifo_cout_drain_out_V_V_din_pass_1_out;
  end
  assign cout_drain_IO_L1_out_wrapper542_U0_fifo_cout_drain_out_V_V_din_pass_1_in = cout_drain_IO_L1_out_wrapper542_U0_fifo_cout_drain_out_V_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_cout_drain_IO_L1_out_10_0_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_cout_drain_IO_L1_out_10_0_V_V_full_n_pass_0_q0 <= fifo_cout_drain_cout_drain_IO_L1_out_10_0_V_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_cout_drain_IO_L1_out_10_0_V_V_full_n_pass_0_in = fifo_cout_drain_cout_drain_IO_L1_out_10_0_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  cout_drain_IO_L1_out_wrapper542_U0_fifo_cout_drain_out_V_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper542_U0_fifo_cout_drain_out_V_V_write_pass_1_q0 <= cout_drain_IO_L1_out_wrapper542_U0_fifo_cout_drain_out_V_V_write_pass_1_out;
  end
  assign cout_drain_IO_L1_out_wrapper542_U0_fifo_cout_drain_out_V_V_write_pass_1_in = cout_drain_IO_L1_out_wrapper542_U0_fifo_cout_drain_out_V_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper219_U0_fifo_cin_out_V_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper219_U0_fifo_cin_out_V_V_din_pass_1_q0 <= PE_wrapper219_U0_fifo_cin_out_V_V_din_pass_1_out;
  end
  assign PE_wrapper219_U0_fifo_cin_out_V_V_din_pass_1_in = PE_wrapper219_U0_fifo_cin_out_V_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_6_9_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_6_9_V_V_full_n_pass_0_q0 <= fifo_cin_PE_6_9_V_V_full_n_pass_0_out;
  end
  assign fifo_cin_PE_6_9_V_V_full_n_pass_0_in = fifo_cin_PE_6_9_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper219_U0_fifo_cin_out_V_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper219_U0_fifo_cin_out_V_V_write_pass_1_q0 <= PE_wrapper219_U0_fifo_cin_out_V_V_write_pass_1_out;
  end
  assign PE_wrapper219_U0_fifo_cin_out_V_V_write_pass_1_in = PE_wrapper219_U0_fifo_cin_out_V_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper172_U0_fifo_cin_out_V_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper172_U0_fifo_cin_out_V_V_din_pass_1_q0 <= PE_wrapper172_U0_fifo_cin_out_V_V_din_pass_1_out;
  end
  assign PE_wrapper172_U0_fifo_cin_out_V_V_din_pass_1_in = PE_wrapper172_U0_fifo_cin_out_V_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_2_10_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_2_10_V_V_full_n_pass_0_q0 <= fifo_cin_PE_2_10_V_V_full_n_pass_0_out;
  end
  assign fifo_cin_PE_2_10_V_V_full_n_pass_0_in = fifo_cin_PE_2_10_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper172_U0_fifo_cin_out_V_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper172_U0_fifo_cin_out_V_V_write_pass_1_q0 <= PE_wrapper172_U0_fifo_cin_out_V_V_write_pass_1_out;
  end
  assign PE_wrapper172_U0_fifo_cin_out_V_V_write_pass_1_in = PE_wrapper172_U0_fifo_cin_out_V_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [255:0] cin_IO_L2_in134_U0_fifo_cin_out_V_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    cin_IO_L2_in134_U0_fifo_cin_out_V_V_din_pass_1_q0 <= cin_IO_L2_in134_U0_fifo_cin_out_V_V_din_pass_1_out;
  end
  assign cin_IO_L2_in134_U0_fifo_cin_out_V_V_din_pass_1_in = cin_IO_L2_in134_U0_fifo_cin_out_V_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_cin_IO_L2_in_11_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_cin_IO_L2_in_11_V_V_full_n_pass_0_q0 <= fifo_cin_cin_IO_L2_in_11_V_V_full_n_pass_0_out;
  end
  assign fifo_cin_cin_IO_L2_in_11_V_V_full_n_pass_0_in = fifo_cin_cin_IO_L2_in_11_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  cin_IO_L2_in134_U0_fifo_cin_out_V_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    cin_IO_L2_in134_U0_fifo_cin_out_V_V_write_pass_1_q0 <= cin_IO_L2_in134_U0_fifo_cin_out_V_V_write_pass_1_out;
  end
  assign cin_IO_L2_in134_U0_fifo_cin_out_V_V_write_pass_1_in = cin_IO_L2_in134_U0_fifo_cin_out_V_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper194_U0_fifo_w_out_V_V_din_pass_2_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper194_U0_fifo_w_out_V_V_din_pass_2_q0 <= PE_wrapper194_U0_fifo_w_out_V_V_din_pass_2_out;
  end
  assign PE_wrapper194_U0_fifo_w_out_V_V_din_pass_2_in = PE_wrapper194_U0_fifo_w_out_V_V_din_pass_2_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_3_9_V_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_3_9_V_V_full_n_pass_1_q0 <= fifo_w_PE_3_9_V_V_full_n_pass_1_out;
  end
  assign fifo_w_PE_3_9_V_V_full_n_pass_1_in = fifo_w_PE_3_9_V_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper194_U0_fifo_w_out_V_V_write_pass_2_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper194_U0_fifo_w_out_V_V_write_pass_2_q0 <= PE_wrapper194_U0_fifo_w_out_V_V_write_pass_2_out;
  end
  assign PE_wrapper194_U0_fifo_w_out_V_V_write_pass_2_in = PE_wrapper194_U0_fifo_w_out_V_V_write_pass_2_q0;
  (* dont_touch = "yes" *) reg [63:0] cout_drain_IO_L1_out_wrapper548_U0_fifo_cout_drain_out_V_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper548_U0_fifo_cout_drain_out_V_V_din_pass_1_q0 <= cout_drain_IO_L1_out_wrapper548_U0_fifo_cout_drain_out_V_V_din_pass_1_out;
  end
  assign cout_drain_IO_L1_out_wrapper548_U0_fifo_cout_drain_out_V_V_din_pass_1_in = cout_drain_IO_L1_out_wrapper548_U0_fifo_cout_drain_out_V_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_cout_drain_IO_L1_out_11_9_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_cout_drain_IO_L1_out_11_9_V_V_full_n_pass_0_q0 <= fifo_cout_drain_cout_drain_IO_L1_out_11_9_V_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_cout_drain_IO_L1_out_11_9_V_V_full_n_pass_0_in = fifo_cout_drain_cout_drain_IO_L1_out_11_9_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  cout_drain_IO_L1_out_wrapper548_U0_fifo_cout_drain_out_V_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper548_U0_fifo_cout_drain_out_V_V_write_pass_1_q0 <= cout_drain_IO_L1_out_wrapper548_U0_fifo_cout_drain_out_V_V_write_pass_1_out;
  end
  assign cout_drain_IO_L1_out_wrapper548_U0_fifo_cout_drain_out_V_V_write_pass_1_in = cout_drain_IO_L1_out_wrapper548_U0_fifo_cout_drain_out_V_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [31:0] PE_wrapper219_U0_fifo_cout_drain_out_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper219_U0_fifo_cout_drain_out_V_din_pass_1_q0 <= PE_wrapper219_U0_fifo_cout_drain_out_V_din_pass_1_out;
  end
  assign PE_wrapper219_U0_fifo_cout_drain_out_V_din_pass_1_in = PE_wrapper219_U0_fifo_cout_drain_out_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_PE_5_9_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_PE_5_9_V_full_n_pass_0_q0 <= fifo_cout_drain_PE_5_9_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_PE_5_9_V_full_n_pass_0_in = fifo_cout_drain_PE_5_9_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper219_U0_fifo_cout_drain_out_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper219_U0_fifo_cout_drain_out_V_write_pass_1_q0 <= PE_wrapper219_U0_fifo_cout_drain_out_V_write_pass_1_out;
  end
  assign PE_wrapper219_U0_fifo_cout_drain_out_V_write_pass_1_in = PE_wrapper219_U0_fifo_cout_drain_out_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [63:0] cout_drain_IO_L1_out_wrapper517_U0_fifo_cout_drain_out_V_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper517_U0_fifo_cout_drain_out_V_V_din_pass_1_q0 <= cout_drain_IO_L1_out_wrapper517_U0_fifo_cout_drain_out_V_V_din_pass_1_out;
  end
  assign cout_drain_IO_L1_out_wrapper517_U0_fifo_cout_drain_out_V_V_din_pass_1_in = cout_drain_IO_L1_out_wrapper517_U0_fifo_cout_drain_out_V_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_cout_drain_IO_L1_out_9_9_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_cout_drain_IO_L1_out_9_9_V_V_full_n_pass_0_q0 <= fifo_cout_drain_cout_drain_IO_L1_out_9_9_V_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_cout_drain_IO_L1_out_9_9_V_V_full_n_pass_0_in = fifo_cout_drain_cout_drain_IO_L1_out_9_9_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  cout_drain_IO_L1_out_wrapper517_U0_fifo_cout_drain_out_V_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper517_U0_fifo_cout_drain_out_V_V_write_pass_1_q0 <= cout_drain_IO_L1_out_wrapper517_U0_fifo_cout_drain_out_V_V_write_pass_1_out;
  end
  assign cout_drain_IO_L1_out_wrapper517_U0_fifo_cout_drain_out_V_V_write_pass_1_in = cout_drain_IO_L1_out_wrapper517_U0_fifo_cout_drain_out_V_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [63:0] cout_drain_IO_L1_out_wrapper533_U0_fifo_cout_drain_out_V_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper533_U0_fifo_cout_drain_out_V_V_din_pass_1_q0 <= cout_drain_IO_L1_out_wrapper533_U0_fifo_cout_drain_out_V_V_din_pass_1_out;
  end
  assign cout_drain_IO_L1_out_wrapper533_U0_fifo_cout_drain_out_V_V_din_pass_1_in = cout_drain_IO_L1_out_wrapper533_U0_fifo_cout_drain_out_V_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_cout_drain_IO_L1_out_10_9_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_cout_drain_IO_L1_out_10_9_V_V_full_n_pass_0_q0 <= fifo_cout_drain_cout_drain_IO_L1_out_10_9_V_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_cout_drain_IO_L1_out_10_9_V_V_full_n_pass_0_in = fifo_cout_drain_cout_drain_IO_L1_out_10_9_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  cout_drain_IO_L1_out_wrapper533_U0_fifo_cout_drain_out_V_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper533_U0_fifo_cout_drain_out_V_V_write_pass_1_q0 <= cout_drain_IO_L1_out_wrapper533_U0_fifo_cout_drain_out_V_V_write_pass_1_out;
  end
  assign cout_drain_IO_L1_out_wrapper533_U0_fifo_cout_drain_out_V_V_write_pass_1_in = cout_drain_IO_L1_out_wrapper533_U0_fifo_cout_drain_out_V_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [63:0] cout_drain_IO_L1_out_wrapper535_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper535_U0_fifo_cout_drain_out_V_V_din_pass_0_q0 <= cout_drain_IO_L1_out_wrapper535_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper535_U0_fifo_cout_drain_out_V_V_din_pass_0_in = cout_drain_IO_L1_out_wrapper535_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  cout_drain_IO_L1_out_wrapper535_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper535_U0_fifo_cout_drain_out_V_V_write_pass_0_q0 <= cout_drain_IO_L1_out_wrapper535_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper535_U0_fifo_cout_drain_out_V_V_write_pass_0_in = cout_drain_IO_L1_out_wrapper535_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_5_10_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_5_10_V_V_full_n_pass_0_q0 <= fifo_w_PE_5_10_V_V_full_n_pass_0_out;
  end
  assign fifo_w_PE_5_10_V_V_full_n_pass_0_in = fifo_w_PE_5_10_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg [63:0] cout_drain_IO_L1_out_wrapper537_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper537_U0_fifo_cout_drain_out_V_V_din_pass_0_q0 <= cout_drain_IO_L1_out_wrapper537_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper537_U0_fifo_cout_drain_out_V_V_din_pass_0_in = cout_drain_IO_L1_out_wrapper537_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  cout_drain_IO_L1_out_wrapper537_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper537_U0_fifo_cout_drain_out_V_V_write_pass_0_q0 <= cout_drain_IO_L1_out_wrapper537_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper537_U0_fifo_cout_drain_out_V_V_write_pass_0_in = cout_drain_IO_L1_out_wrapper537_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_2_9_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_2_9_V_V_full_n_pass_0_q0 <= fifo_cin_PE_2_9_V_V_full_n_pass_0_out;
  end
  assign fifo_cin_PE_2_9_V_V_full_n_pass_0_in = fifo_cin_PE_2_9_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_1_11_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_1_11_V_V_full_n_pass_0_q0 <= fifo_w_PE_1_11_V_V_full_n_pass_0_out;
  end
  assign fifo_w_PE_1_11_V_V_full_n_pass_0_in = fifo_w_PE_1_11_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_cout_drain_IO_L1_out_11_6_V_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_cout_drain_IO_L1_out_11_6_V_V_full_n_pass_1_q0 <= fifo_cout_drain_cout_drain_IO_L1_out_11_6_V_V_full_n_pass_1_out;
  end
  assign fifo_cout_drain_cout_drain_IO_L1_out_11_6_V_V_full_n_pass_1_in = fifo_cout_drain_cout_drain_IO_L1_out_11_6_V_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg [63:0] cout_drain_IO_L1_out_wrapper555_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper555_U0_fifo_cout_drain_out_V_V_din_pass_0_q0 <= cout_drain_IO_L1_out_wrapper555_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper555_U0_fifo_cout_drain_out_V_V_din_pass_0_in = cout_drain_IO_L1_out_wrapper555_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  cout_drain_IO_L1_out_wrapper555_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper555_U0_fifo_cout_drain_out_V_V_write_pass_0_q0 <= cout_drain_IO_L1_out_wrapper555_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper555_U0_fifo_cout_drain_out_V_V_write_pass_0_in = cout_drain_IO_L1_out_wrapper555_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_4_10_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_4_10_V_V_full_n_pass_0_q0 <= fifo_cin_PE_4_10_V_V_full_n_pass_0_out;
  end
  assign fifo_cin_PE_4_10_V_V_full_n_pass_0_in = fifo_cin_PE_4_10_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_cout_drain_IO_L1_out_10_3_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_cout_drain_IO_L1_out_10_3_V_V_full_n_pass_0_q0 <= fifo_cout_drain_cout_drain_IO_L1_out_10_3_V_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_cout_drain_IO_L1_out_10_3_V_V_full_n_pass_0_in = fifo_cout_drain_cout_drain_IO_L1_out_10_3_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper244_U0_fifo_cin_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper244_U0_fifo_cin_out_V_V_din_pass_0_q0 <= PE_wrapper244_U0_fifo_cin_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper244_U0_fifo_cin_out_V_V_din_pass_0_in = PE_wrapper244_U0_fifo_cin_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper244_U0_fifo_cin_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper244_U0_fifo_cin_out_V_V_write_pass_0_q0 <= PE_wrapper244_U0_fifo_cin_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper244_U0_fifo_cin_out_V_V_write_pass_0_in = PE_wrapper244_U0_fifo_cin_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_6_10_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_6_10_V_V_full_n_pass_0_q0 <= fifo_w_PE_6_10_V_V_full_n_pass_0_out;
  end
  assign fifo_w_PE_6_10_V_V_full_n_pass_0_in = fifo_w_PE_6_10_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper173_U0_fifo_w_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper173_U0_fifo_w_out_V_V_din_pass_0_q0 <= PE_wrapper173_U0_fifo_w_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper173_U0_fifo_w_out_V_V_din_pass_0_in = PE_wrapper173_U0_fifo_w_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper173_U0_fifo_w_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper173_U0_fifo_w_out_V_V_write_pass_0_q0 <= PE_wrapper173_U0_fifo_w_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper173_U0_fifo_w_out_V_V_write_pass_0_in = PE_wrapper173_U0_fifo_w_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_PE_6_9_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_PE_6_9_V_full_n_pass_0_q0 <= fifo_cout_drain_PE_6_9_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_PE_6_9_V_full_n_pass_0_in = fifo_cout_drain_PE_6_9_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_4_10_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_4_10_V_V_full_n_pass_0_q0 <= fifo_w_PE_4_10_V_V_full_n_pass_0_out;
  end
  assign fifo_w_PE_4_10_V_V_full_n_pass_0_in = fifo_w_PE_4_10_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_PE_5_11_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_PE_5_11_V_full_n_pass_0_q0 <= fifo_cout_drain_PE_5_11_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_PE_5_11_V_full_n_pass_0_in = fifo_cout_drain_PE_5_11_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg [31:0] PE_wrapper183_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper183_U0_fifo_cout_drain_out_V_din_pass_0_q0 <= PE_wrapper183_U0_fifo_cout_drain_out_V_din_pass_0_out;
  end
  assign PE_wrapper183_U0_fifo_cout_drain_out_V_din_pass_0_in = PE_wrapper183_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper183_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper183_U0_fifo_cout_drain_out_V_write_pass_0_q0 <= PE_wrapper183_U0_fifo_cout_drain_out_V_write_pass_0_out;
  end
  assign PE_wrapper183_U0_fifo_cout_drain_out_V_write_pass_0_in = PE_wrapper183_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_1_11_V_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_1_11_V_V_full_n_pass_1_q0 <= fifo_cin_PE_1_11_V_V_full_n_pass_1_out;
  end
  assign fifo_cin_PE_1_11_V_V_full_n_pass_1_in = fifo_cin_PE_1_11_V_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg [31:0] PE_wrapper232_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper232_U0_fifo_cout_drain_out_V_din_pass_0_q0 <= PE_wrapper232_U0_fifo_cout_drain_out_V_din_pass_0_out;
  end
  assign PE_wrapper232_U0_fifo_cout_drain_out_V_din_pass_0_in = PE_wrapper232_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper232_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper232_U0_fifo_cout_drain_out_V_write_pass_0_q0 <= PE_wrapper232_U0_fifo_cout_drain_out_V_write_pass_0_out;
  end
  assign PE_wrapper232_U0_fifo_cout_drain_out_V_write_pass_0_in = PE_wrapper232_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  cout_V_c_full_n_pass_5_q0;
  always @ (posedge ap_clk) begin
    cout_V_c_full_n_pass_5_q0 <= cout_V_c_full_n_pass_5_out;
  end
  assign cout_V_c_full_n_pass_5_in = cout_V_c_full_n_pass_5_q0;
  (* dont_touch = "yes" *) reg [63:0] cout_drain_IO_L1_out_wrapper540_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper540_U0_fifo_cout_drain_out_V_V_din_pass_0_q0 <= cout_drain_IO_L1_out_wrapper540_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper540_U0_fifo_cout_drain_out_V_V_din_pass_0_in = cout_drain_IO_L1_out_wrapper540_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  cout_drain_IO_L1_out_wrapper540_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper540_U0_fifo_cout_drain_out_V_V_write_pass_0_q0 <= cout_drain_IO_L1_out_wrapper540_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper540_U0_fifo_cout_drain_out_V_V_write_pass_0_in = cout_drain_IO_L1_out_wrapper540_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [63:0] cout_drain_IO_L1_out_wrapper552_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper552_U0_fifo_cout_drain_out_V_V_din_pass_0_q0 <= cout_drain_IO_L1_out_wrapper552_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper552_U0_fifo_cout_drain_out_V_V_din_pass_0_in = cout_drain_IO_L1_out_wrapper552_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  cout_drain_IO_L1_out_wrapper552_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper552_U0_fifo_cout_drain_out_V_V_write_pass_0_q0 <= cout_drain_IO_L1_out_wrapper552_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper552_U0_fifo_cout_drain_out_V_V_write_pass_0_in = cout_drain_IO_L1_out_wrapper552_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_7_10_V_V_full_n_pass_3_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_7_10_V_V_full_n_pass_3_q0 <= fifo_w_PE_7_10_V_V_full_n_pass_3_out;
  end
  assign fifo_w_PE_7_10_V_V_full_n_pass_3_in = fifo_w_PE_7_10_V_V_full_n_pass_3_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_PE_7_9_V_full_n_pass_3_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_PE_7_9_V_full_n_pass_3_q0 <= fifo_cout_drain_PE_7_9_V_full_n_pass_3_out;
  end
  assign fifo_cout_drain_PE_7_9_V_full_n_pass_3_in = fifo_cout_drain_PE_7_9_V_full_n_pass_3_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_PE_2_10_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_PE_2_10_V_full_n_pass_0_q0 <= fifo_cout_drain_PE_2_10_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_PE_2_10_V_full_n_pass_0_in = fifo_cout_drain_PE_2_10_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_8_9_V_V_full_n_pass_3_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_8_9_V_V_full_n_pass_3_q0 <= fifo_cin_PE_8_9_V_V_full_n_pass_3_out;
  end
  assign fifo_cin_PE_8_9_V_V_full_n_pass_3_in = fifo_cin_PE_8_9_V_V_full_n_pass_3_q0;
  (* dont_touch = "yes" *) reg [31:0] PE_wrapper255_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper255_U0_fifo_cout_drain_out_V_din_pass_0_q0 <= PE_wrapper255_U0_fifo_cout_drain_out_V_din_pass_0_out;
  end
  assign PE_wrapper255_U0_fifo_cout_drain_out_V_din_pass_0_in = PE_wrapper255_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper255_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper255_U0_fifo_cout_drain_out_V_write_pass_0_q0 <= PE_wrapper255_U0_fifo_cout_drain_out_V_write_pass_0_out;
  end
  assign PE_wrapper255_U0_fifo_cout_drain_out_V_write_pass_0_in = PE_wrapper255_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_PE_2_11_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_PE_2_11_V_full_n_pass_1_q0 <= fifo_cout_drain_PE_2_11_V_full_n_pass_1_out;
  end
  assign fifo_cout_drain_PE_2_11_V_full_n_pass_1_in = fifo_cout_drain_PE_2_11_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_cout_drain_IO_L1_out_9_8_V_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_cout_drain_IO_L1_out_9_8_V_V_full_n_pass_1_q0 <= fifo_cout_drain_cout_drain_IO_L1_out_9_8_V_V_full_n_pass_1_out;
  end
  assign fifo_cout_drain_cout_drain_IO_L1_out_9_8_V_V_full_n_pass_1_in = fifo_cout_drain_cout_drain_IO_L1_out_9_8_V_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper255_U0_fifo_cin_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper255_U0_fifo_cin_out_V_V_din_pass_0_q0 <= PE_wrapper255_U0_fifo_cin_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper255_U0_fifo_cin_out_V_V_din_pass_0_in = PE_wrapper255_U0_fifo_cin_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper255_U0_fifo_cin_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper255_U0_fifo_cin_out_V_V_write_pass_0_q0 <= PE_wrapper255_U0_fifo_cin_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper255_U0_fifo_cin_out_V_V_write_pass_0_in = PE_wrapper255_U0_fifo_cin_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper244_U0_fifo_w_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper244_U0_fifo_w_out_V_V_din_pass_0_q0 <= PE_wrapper244_U0_fifo_w_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper244_U0_fifo_w_out_V_V_din_pass_0_in = PE_wrapper244_U0_fifo_w_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper244_U0_fifo_w_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper244_U0_fifo_w_out_V_V_write_pass_0_q0 <= PE_wrapper244_U0_fifo_w_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper244_U0_fifo_w_out_V_V_write_pass_0_in = PE_wrapper244_U0_fifo_w_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [31:0] PE_wrapper173_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper173_U0_fifo_cout_drain_out_V_din_pass_0_q0 <= PE_wrapper173_U0_fifo_cout_drain_out_V_din_pass_0_out;
  end
  assign PE_wrapper173_U0_fifo_cout_drain_out_V_din_pass_0_in = PE_wrapper173_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper173_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper173_U0_fifo_cout_drain_out_V_write_pass_0_q0 <= PE_wrapper173_U0_fifo_cout_drain_out_V_write_pass_0_out;
  end
  assign PE_wrapper173_U0_fifo_cout_drain_out_V_write_pass_0_in = PE_wrapper173_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_8_9_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_8_9_V_V_full_n_pass_0_q0 <= fifo_w_PE_8_9_V_V_full_n_pass_0_out;
  end
  assign fifo_w_PE_8_9_V_V_full_n_pass_0_in = fifo_w_PE_8_9_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg [31:0] PE_wrapper208_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper208_U0_fifo_cout_drain_out_V_din_pass_0_q0 <= PE_wrapper208_U0_fifo_cout_drain_out_V_din_pass_0_out;
  end
  assign PE_wrapper208_U0_fifo_cout_drain_out_V_din_pass_0_in = PE_wrapper208_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper208_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper208_U0_fifo_cout_drain_out_V_write_pass_0_q0 <= PE_wrapper208_U0_fifo_cout_drain_out_V_write_pass_0_out;
  end
  assign PE_wrapper208_U0_fifo_cout_drain_out_V_write_pass_0_in = PE_wrapper208_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_cout_drain_IO_L1_out_10_6_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_cout_drain_IO_L1_out_10_6_V_V_full_n_pass_0_q0 <= fifo_cout_drain_cout_drain_IO_L1_out_10_6_V_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_cout_drain_IO_L1_out_10_6_V_V_full_n_pass_0_in = fifo_cout_drain_cout_drain_IO_L1_out_10_6_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_2_9_V_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_2_9_V_V_full_n_pass_1_q0 <= fifo_w_PE_2_9_V_V_full_n_pass_1_out;
  end
  assign fifo_w_PE_2_9_V_V_full_n_pass_1_in = fifo_w_PE_2_9_V_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper220_U0_fifo_w_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper220_U0_fifo_w_out_V_V_din_pass_0_q0 <= PE_wrapper220_U0_fifo_w_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper220_U0_fifo_w_out_V_V_din_pass_0_in = PE_wrapper220_U0_fifo_w_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper220_U0_fifo_w_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper220_U0_fifo_w_out_V_V_write_pass_0_q0 <= PE_wrapper220_U0_fifo_w_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper220_U0_fifo_w_out_V_V_write_pass_0_in = PE_wrapper220_U0_fifo_w_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper255_U0_fifo_w_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper255_U0_fifo_w_out_V_V_din_pass_0_q0 <= PE_wrapper255_U0_fifo_w_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper255_U0_fifo_w_out_V_V_din_pass_0_in = PE_wrapper255_U0_fifo_w_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper255_U0_fifo_w_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper255_U0_fifo_w_out_V_V_write_pass_0_q0 <= PE_wrapper255_U0_fifo_w_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper255_U0_fifo_w_out_V_V_write_pass_0_in = PE_wrapper255_U0_fifo_w_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_cout_drain_IO_L1_out_10_8_V_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_cout_drain_IO_L1_out_10_8_V_V_full_n_pass_1_q0 <= fifo_cout_drain_cout_drain_IO_L1_out_10_8_V_V_full_n_pass_1_out;
  end
  assign fifo_cout_drain_cout_drain_IO_L1_out_10_8_V_V_full_n_pass_1_in = fifo_cout_drain_cout_drain_IO_L1_out_10_8_V_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg [63:0] cout_drain_IO_L1_out_wrapper520_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper520_U0_fifo_cout_drain_out_V_V_din_pass_0_q0 <= cout_drain_IO_L1_out_wrapper520_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper520_U0_fifo_cout_drain_out_V_V_din_pass_0_in = cout_drain_IO_L1_out_wrapper520_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  cout_drain_IO_L1_out_wrapper520_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper520_U0_fifo_cout_drain_out_V_V_write_pass_0_q0 <= cout_drain_IO_L1_out_wrapper520_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper520_U0_fifo_cout_drain_out_V_V_write_pass_0_in = cout_drain_IO_L1_out_wrapper520_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_cout_drain_IO_L3_out_serialize_V_V_full_n_pass_2_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_cout_drain_IO_L3_out_serialize_V_V_full_n_pass_2_q0 <= fifo_cout_drain_cout_drain_IO_L3_out_serialize_V_V_full_n_pass_2_out;
  end
  assign fifo_cout_drain_cout_drain_IO_L3_out_serialize_V_V_full_n_pass_2_in = fifo_cout_drain_cout_drain_IO_L3_out_serialize_V_V_full_n_pass_2_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper173_U0_fifo_cin_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper173_U0_fifo_cin_out_V_V_din_pass_0_q0 <= PE_wrapper173_U0_fifo_cin_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper173_U0_fifo_cin_out_V_V_din_pass_0_in = PE_wrapper173_U0_fifo_cin_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper173_U0_fifo_cin_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper173_U0_fifo_cin_out_V_V_write_pass_0_q0 <= PE_wrapper173_U0_fifo_cin_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper173_U0_fifo_cin_out_V_V_write_pass_0_in = PE_wrapper173_U0_fifo_cin_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper232_U0_fifo_w_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper232_U0_fifo_w_out_V_V_din_pass_0_q0 <= PE_wrapper232_U0_fifo_w_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper232_U0_fifo_w_out_V_V_din_pass_0_in = PE_wrapper232_U0_fifo_w_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper232_U0_fifo_w_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper232_U0_fifo_w_out_V_V_write_pass_0_q0 <= PE_wrapper232_U0_fifo_w_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper232_U0_fifo_w_out_V_V_write_pass_0_in = PE_wrapper232_U0_fifo_w_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper183_U0_fifo_w_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper183_U0_fifo_w_out_V_V_din_pass_0_q0 <= PE_wrapper183_U0_fifo_w_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper183_U0_fifo_w_out_V_V_din_pass_0_in = PE_wrapper183_U0_fifo_w_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper183_U0_fifo_w_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper183_U0_fifo_w_out_V_V_write_pass_0_q0 <= PE_wrapper183_U0_fifo_w_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper183_U0_fifo_w_out_V_V_write_pass_0_in = PE_wrapper183_U0_fifo_w_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_5_12_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_5_12_V_V_full_n_pass_0_q0 <= fifo_w_PE_5_12_V_V_full_n_pass_0_out;
  end
  assign fifo_w_PE_5_12_V_V_full_n_pass_0_in = fifo_w_PE_5_12_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper208_U0_fifo_w_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper208_U0_fifo_w_out_V_V_din_pass_0_q0 <= PE_wrapper208_U0_fifo_w_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper208_U0_fifo_w_out_V_V_din_pass_0_in = PE_wrapper208_U0_fifo_w_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper208_U0_fifo_w_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper208_U0_fifo_w_out_V_V_write_pass_0_q0 <= PE_wrapper208_U0_fifo_w_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper208_U0_fifo_w_out_V_V_write_pass_0_in = PE_wrapper208_U0_fifo_w_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_PE_3_11_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_PE_3_11_V_full_n_pass_1_q0 <= fifo_cout_drain_PE_3_11_V_full_n_pass_1_out;
  end
  assign fifo_cout_drain_PE_3_11_V_full_n_pass_1_in = fifo_cout_drain_PE_3_11_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper183_U0_fifo_cin_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper183_U0_fifo_cin_out_V_V_din_pass_0_q0 <= PE_wrapper183_U0_fifo_cin_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper183_U0_fifo_cin_out_V_V_din_pass_0_in = PE_wrapper183_U0_fifo_cin_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper183_U0_fifo_cin_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper183_U0_fifo_cin_out_V_V_write_pass_0_q0 <= PE_wrapper183_U0_fifo_cin_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper183_U0_fifo_cin_out_V_V_write_pass_0_in = PE_wrapper183_U0_fifo_cin_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_cout_drain_IO_L1_out_11_4_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_cout_drain_IO_L1_out_11_4_V_V_full_n_pass_0_q0 <= fifo_cout_drain_cout_drain_IO_L1_out_11_4_V_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_cout_drain_IO_L1_out_11_4_V_V_full_n_pass_0_in = fifo_cout_drain_cout_drain_IO_L1_out_11_4_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  ap_done_Boundary_X4Y12_To_X6Y12_q0;
  always @ (posedge ap_clk) begin
    ap_done_Boundary_X4Y12_To_X6Y12_q0 <= ap_done_Boundary_X4Y12_To_X6Y12_out;
  end
  assign ap_done_Boundary_X4Y12_To_X6Y12_in = ap_done_Boundary_X4Y12_To_X6Y12_q0;
  (* dont_touch = "yes" *) reg  ap_start_Boundary_X4Y14_To_X6Y14_q0;
  always @ (posedge ap_clk) begin
    ap_start_Boundary_X4Y14_To_X6Y14_q0 <= ap_start_Boundary_X4Y14_To_X6Y14_out;
  end
  assign ap_start_Boundary_X4Y14_To_X6Y14_in = ap_start_Boundary_X4Y14_To_X6Y14_q0;
  (* dont_touch = "yes" *) reg  ap_rst_n_Boundary_X4Y14_To_X6Y14_q0;
  always @ (posedge ap_clk) begin
    ap_rst_n_Boundary_X4Y14_To_X6Y14_q0 <= ap_rst_n_Boundary_X4Y14_To_X6Y14_out;
  end
  assign ap_rst_n_Boundary_X4Y14_To_X6Y14_in = ap_rst_n_Boundary_X4Y14_To_X6Y14_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper260_U0_fifo_cin_out_V_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper260_U0_fifo_cin_out_V_V_din_pass_1_q0 <= PE_wrapper260_U0_fifo_cin_out_V_V_din_pass_1_out;
  end
  assign PE_wrapper260_U0_fifo_cin_out_V_V_din_pass_1_in = PE_wrapper260_U0_fifo_cin_out_V_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_10_2_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_10_2_V_V_full_n_pass_0_q0 <= fifo_cin_PE_10_2_V_V_full_n_pass_0_out;
  end
  assign fifo_cin_PE_10_2_V_V_full_n_pass_0_in = fifo_cin_PE_10_2_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper260_U0_fifo_cin_out_V_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper260_U0_fifo_cin_out_V_V_write_pass_1_q0 <= PE_wrapper260_U0_fifo_cin_out_V_V_write_pass_1_out;
  end
  assign PE_wrapper260_U0_fifo_cin_out_V_V_write_pass_1_in = PE_wrapper260_U0_fifo_cin_out_V_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper261_U0_fifo_w_out_V_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper261_U0_fifo_w_out_V_V_din_pass_1_q0 <= PE_wrapper261_U0_fifo_w_out_V_V_din_pass_1_out;
  end
  assign PE_wrapper261_U0_fifo_w_out_V_V_din_pass_1_in = PE_wrapper261_U0_fifo_w_out_V_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_9_4_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_9_4_V_V_full_n_pass_0_q0 <= fifo_w_PE_9_4_V_V_full_n_pass_0_out;
  end
  assign fifo_w_PE_9_4_V_V_full_n_pass_0_in = fifo_w_PE_9_4_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper261_U0_fifo_w_out_V_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper261_U0_fifo_w_out_V_V_write_pass_1_q0 <= PE_wrapper261_U0_fifo_w_out_V_V_write_pass_1_out;
  end
  assign PE_wrapper261_U0_fifo_w_out_V_V_write_pass_1_in = PE_wrapper261_U0_fifo_w_out_V_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [255:0] w_IO_L2_in144_U0_fifo_w_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    w_IO_L2_in144_U0_fifo_w_out_V_V_din_pass_0_q0 <= w_IO_L2_in144_U0_fifo_w_out_V_V_din_pass_0_out;
  end
  assign w_IO_L2_in144_U0_fifo_w_out_V_V_din_pass_0_in = w_IO_L2_in144_U0_fifo_w_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  w_IO_L2_in144_U0_fifo_w_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    w_IO_L2_in144_U0_fifo_w_out_V_V_write_pass_0_q0 <= w_IO_L2_in144_U0_fifo_w_out_V_V_write_pass_0_out;
  end
  assign w_IO_L2_in144_U0_fifo_w_out_V_V_write_pass_0_in = w_IO_L2_in144_U0_fifo_w_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [31:0] PE_wrapper271_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper271_U0_fifo_cout_drain_out_V_din_pass_0_q0 <= PE_wrapper271_U0_fifo_cout_drain_out_V_din_pass_0_out;
  end
  assign PE_wrapper271_U0_fifo_cout_drain_out_V_din_pass_0_in = PE_wrapper271_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper271_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper271_U0_fifo_cout_drain_out_V_write_pass_0_q0 <= PE_wrapper271_U0_fifo_cout_drain_out_V_write_pass_0_out;
  end
  assign PE_wrapper271_U0_fifo_cout_drain_out_V_write_pass_0_in = PE_wrapper271_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_cout_drain_IO_L1_out_0_10_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_cout_drain_IO_L1_out_0_10_V_V_full_n_pass_0_q0 <= fifo_cout_drain_cout_drain_IO_L1_out_0_10_V_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_cout_drain_IO_L1_out_0_10_V_V_full_n_pass_0_in = fifo_cout_drain_cout_drain_IO_L1_out_0_10_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg [31:0] PE_wrapper247_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper247_U0_fifo_cout_drain_out_V_din_pass_0_q0 <= PE_wrapper247_U0_fifo_cout_drain_out_V_din_pass_0_out;
  end
  assign PE_wrapper247_U0_fifo_cout_drain_out_V_din_pass_0_in = PE_wrapper247_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper247_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper247_U0_fifo_cout_drain_out_V_write_pass_0_q0 <= PE_wrapper247_U0_fifo_cout_drain_out_V_write_pass_0_out;
  end
  assign PE_wrapper247_U0_fifo_cout_drain_out_V_write_pass_0_in = PE_wrapper247_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [31:0] PE_wrapper259_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper259_U0_fifo_cout_drain_out_V_din_pass_0_q0 <= PE_wrapper259_U0_fifo_cout_drain_out_V_din_pass_0_out;
  end
  assign PE_wrapper259_U0_fifo_cout_drain_out_V_din_pass_0_in = PE_wrapper259_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper259_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper259_U0_fifo_cout_drain_out_V_write_pass_0_q0 <= PE_wrapper259_U0_fifo_cout_drain_out_V_write_pass_0_out;
  end
  assign PE_wrapper259_U0_fifo_cout_drain_out_V_write_pass_0_in = PE_wrapper259_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_8_0_V_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_8_0_V_V_full_n_pass_1_q0 <= fifo_cin_PE_8_0_V_V_full_n_pass_1_out;
  end
  assign fifo_cin_PE_8_0_V_V_full_n_pass_1_in = fifo_cin_PE_8_0_V_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper258_U0_fifo_cin_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper258_U0_fifo_cin_out_V_V_din_pass_0_q0 <= PE_wrapper258_U0_fifo_cin_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper258_U0_fifo_cin_out_V_V_din_pass_0_in = PE_wrapper258_U0_fifo_cin_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper258_U0_fifo_cin_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper258_U0_fifo_cin_out_V_V_write_pass_0_q0 <= PE_wrapper258_U0_fifo_cin_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper258_U0_fifo_cin_out_V_V_write_pass_0_in = PE_wrapper258_U0_fifo_cin_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [63:0] cout_drain_IO_L1_out_wrapper374_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper374_U0_fifo_cout_drain_out_V_V_din_pass_0_q0 <= cout_drain_IO_L1_out_wrapper374_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper374_U0_fifo_cout_drain_out_V_V_din_pass_0_in = cout_drain_IO_L1_out_wrapper374_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  cout_drain_IO_L1_out_wrapper374_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper374_U0_fifo_cout_drain_out_V_V_write_pass_0_q0 <= cout_drain_IO_L1_out_wrapper374_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper374_U0_fifo_cout_drain_out_V_V_write_pass_0_in = cout_drain_IO_L1_out_wrapper374_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_8_1_V_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_8_1_V_V_full_n_pass_1_q0 <= fifo_cin_PE_8_1_V_V_full_n_pass_1_out;
  end
  assign fifo_cin_PE_8_1_V_V_full_n_pass_1_in = fifo_cin_PE_8_1_V_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper247_U0_fifo_w_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper247_U0_fifo_w_out_V_V_din_pass_0_q0 <= PE_wrapper247_U0_fifo_w_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper247_U0_fifo_w_out_V_V_din_pass_0_in = PE_wrapper247_U0_fifo_w_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper247_U0_fifo_w_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper247_U0_fifo_w_out_V_V_write_pass_0_q0 <= PE_wrapper247_U0_fifo_w_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper247_U0_fifo_w_out_V_V_write_pass_0_in = PE_wrapper247_U0_fifo_w_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_w_w_IO_L2_in_8_V_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_w_w_IO_L2_in_8_V_V_full_n_pass_1_q0 <= fifo_w_w_IO_L2_in_8_V_V_full_n_pass_1_out;
  end
  assign fifo_w_w_IO_L2_in_8_V_V_full_n_pass_1_in = fifo_w_w_IO_L2_in_8_V_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper271_U0_fifo_cin_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper271_U0_fifo_cin_out_V_V_din_pass_0_q0 <= PE_wrapper271_U0_fifo_cin_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper271_U0_fifo_cin_out_V_V_din_pass_0_in = PE_wrapper271_U0_fifo_cin_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper271_U0_fifo_cin_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper271_U0_fifo_cin_out_V_V_write_pass_0_q0 <= PE_wrapper271_U0_fifo_cin_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper271_U0_fifo_cin_out_V_V_write_pass_0_in = PE_wrapper271_U0_fifo_cin_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_10_1_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_10_1_V_V_full_n_pass_0_q0 <= fifo_w_PE_10_1_V_V_full_n_pass_0_out;
  end
  assign fifo_w_PE_10_1_V_V_full_n_pass_0_in = fifo_w_PE_10_1_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper259_U0_fifo_w_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper259_U0_fifo_w_out_V_V_din_pass_0_q0 <= PE_wrapper259_U0_fifo_w_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper259_U0_fifo_w_out_V_V_din_pass_0_in = PE_wrapper259_U0_fifo_w_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper259_U0_fifo_w_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper259_U0_fifo_w_out_V_V_write_pass_0_q0 <= PE_wrapper259_U0_fifo_w_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper259_U0_fifo_w_out_V_V_write_pass_0_in = PE_wrapper259_U0_fifo_w_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper271_U0_fifo_w_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper271_U0_fifo_w_out_V_V_din_pass_0_q0 <= PE_wrapper271_U0_fifo_w_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper271_U0_fifo_w_out_V_V_din_pass_0_in = PE_wrapper271_U0_fifo_w_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper271_U0_fifo_w_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper271_U0_fifo_w_out_V_V_write_pass_0_q0 <= PE_wrapper271_U0_fifo_w_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper271_U0_fifo_w_out_V_V_write_pass_0_in = PE_wrapper271_U0_fifo_w_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  ap_done_Boundary_X2Y0_To_X2Y2_q0;
  always @ (posedge ap_clk) begin
    ap_done_Boundary_X2Y0_To_X2Y2_q0 <= ap_done_Boundary_X2Y0_To_X2Y2_out;
  end
  assign ap_done_Boundary_X2Y0_To_X2Y2_in = ap_done_Boundary_X2Y0_To_X2Y2_q0;
  (* dont_touch = "yes" *) reg  ap_start_Boundary_X0Y2_To_X2Y2_q0;
  always @ (posedge ap_clk) begin
    ap_start_Boundary_X0Y2_To_X2Y2_q0 <= ap_start_Boundary_X0Y2_To_X2Y2_out;
  end
  assign ap_start_Boundary_X0Y2_To_X2Y2_in = ap_start_Boundary_X0Y2_To_X2Y2_q0;
  (* dont_touch = "yes" *) reg  ap_rst_n_Boundary_X0Y2_To_X2Y2_q0;
  always @ (posedge ap_clk) begin
    ap_rst_n_Boundary_X0Y2_To_X2Y2_q0 <= ap_rst_n_Boundary_X0Y2_To_X2Y2_out;
  end
  assign ap_rst_n_Boundary_X0Y2_To_X2Y2_in = ap_rst_n_Boundary_X0Y2_To_X2Y2_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper234_U0_fifo_cin_out_V_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper234_U0_fifo_cin_out_V_V_din_pass_1_q0 <= PE_wrapper234_U0_fifo_cin_out_V_V_din_pass_1_out;
  end
  assign PE_wrapper234_U0_fifo_cin_out_V_V_din_pass_1_in = PE_wrapper234_U0_fifo_cin_out_V_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_8_0_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_8_0_V_V_full_n_pass_0_q0 <= fifo_cin_PE_8_0_V_V_full_n_pass_0_out;
  end
  assign fifo_cin_PE_8_0_V_V_full_n_pass_0_in = fifo_cin_PE_8_0_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper234_U0_fifo_cin_out_V_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper234_U0_fifo_cin_out_V_V_write_pass_1_q0 <= PE_wrapper234_U0_fifo_cin_out_V_V_write_pass_1_out;
  end
  assign PE_wrapper234_U0_fifo_cin_out_V_V_write_pass_1_in = PE_wrapper234_U0_fifo_cin_out_V_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper235_U0_fifo_cin_out_V_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper235_U0_fifo_cin_out_V_V_din_pass_1_q0 <= PE_wrapper235_U0_fifo_cin_out_V_V_din_pass_1_out;
  end
  assign PE_wrapper235_U0_fifo_cin_out_V_V_din_pass_1_in = PE_wrapper235_U0_fifo_cin_out_V_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_8_1_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_8_1_V_V_full_n_pass_0_q0 <= fifo_cin_PE_8_1_V_V_full_n_pass_0_out;
  end
  assign fifo_cin_PE_8_1_V_V_full_n_pass_0_in = fifo_cin_PE_8_1_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper235_U0_fifo_cin_out_V_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper235_U0_fifo_cin_out_V_V_write_pass_1_q0 <= PE_wrapper235_U0_fifo_cin_out_V_V_write_pass_1_out;
  end
  assign PE_wrapper235_U0_fifo_cin_out_V_V_write_pass_1_in = PE_wrapper235_U0_fifo_cin_out_V_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [255:0] w_IO_L2_in142_U0_fifo_w_out_V_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    w_IO_L2_in142_U0_fifo_w_out_V_V_din_pass_1_q0 <= w_IO_L2_in142_U0_fifo_w_out_V_V_din_pass_1_out;
  end
  assign w_IO_L2_in142_U0_fifo_w_out_V_V_din_pass_1_in = w_IO_L2_in142_U0_fifo_w_out_V_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_w_w_IO_L2_in_8_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_w_IO_L2_in_8_V_V_full_n_pass_0_q0 <= fifo_w_w_IO_L2_in_8_V_V_full_n_pass_0_out;
  end
  assign fifo_w_w_IO_L2_in_8_V_V_full_n_pass_0_in = fifo_w_w_IO_L2_in_8_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  w_IO_L2_in142_U0_fifo_w_out_V_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    w_IO_L2_in142_U0_fifo_w_out_V_V_write_pass_1_q0 <= w_IO_L2_in142_U0_fifo_w_out_V_V_write_pass_1_out;
  end
  assign w_IO_L2_in142_U0_fifo_w_out_V_V_write_pass_1_in = w_IO_L2_in142_U0_fifo_w_out_V_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper261_U0_fifo_w_out_V_V_din_pass_2_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper261_U0_fifo_w_out_V_V_din_pass_2_q0 <= PE_wrapper261_U0_fifo_w_out_V_V_din_pass_2_out;
  end
  assign PE_wrapper261_U0_fifo_w_out_V_V_din_pass_2_in = PE_wrapper261_U0_fifo_w_out_V_V_din_pass_2_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_9_4_V_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_9_4_V_V_full_n_pass_1_q0 <= fifo_w_PE_9_4_V_V_full_n_pass_1_out;
  end
  assign fifo_w_PE_9_4_V_V_full_n_pass_1_in = fifo_w_PE_9_4_V_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper261_U0_fifo_w_out_V_V_write_pass_2_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper261_U0_fifo_w_out_V_V_write_pass_2_q0 <= PE_wrapper261_U0_fifo_w_out_V_V_write_pass_2_out;
  end
  assign PE_wrapper261_U0_fifo_w_out_V_V_write_pass_2_in = PE_wrapper261_U0_fifo_w_out_V_V_write_pass_2_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper237_U0_fifo_w_out_V_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper237_U0_fifo_w_out_V_V_din_pass_1_q0 <= PE_wrapper237_U0_fifo_w_out_V_V_din_pass_1_out;
  end
  assign PE_wrapper237_U0_fifo_w_out_V_V_din_pass_1_in = PE_wrapper237_U0_fifo_w_out_V_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_7_4_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_7_4_V_V_full_n_pass_0_q0 <= fifo_w_PE_7_4_V_V_full_n_pass_0_out;
  end
  assign fifo_w_PE_7_4_V_V_full_n_pass_0_in = fifo_w_PE_7_4_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper237_U0_fifo_w_out_V_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper237_U0_fifo_w_out_V_V_write_pass_1_q0 <= PE_wrapper237_U0_fifo_w_out_V_V_write_pass_1_out;
  end
  assign PE_wrapper237_U0_fifo_w_out_V_V_write_pass_1_in = PE_wrapper237_U0_fifo_w_out_V_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_10_2_V_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_10_2_V_V_full_n_pass_1_q0 <= fifo_cin_PE_10_2_V_V_full_n_pass_1_out;
  end
  assign fifo_cin_PE_10_2_V_V_full_n_pass_1_in = fifo_cin_PE_10_2_V_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_cout_drain_IO_L1_out_2_12_V_V_full_n_pass_2_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_cout_drain_IO_L1_out_2_12_V_V_full_n_pass_2_q0 <= fifo_cout_drain_cout_drain_IO_L1_out_2_12_V_V_full_n_pass_2_out;
  end
  assign fifo_cout_drain_cout_drain_IO_L1_out_2_12_V_V_full_n_pass_2_in = fifo_cout_drain_cout_drain_IO_L1_out_2_12_V_V_full_n_pass_2_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_10_2_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_10_2_V_V_full_n_pass_0_q0 <= fifo_w_PE_10_2_V_V_full_n_pass_0_out;
  end
  assign fifo_w_PE_10_2_V_V_full_n_pass_0_in = fifo_w_PE_10_2_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg [63:0] cout_drain_IO_L1_out_wrapper372_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper372_U0_fifo_cout_drain_out_V_V_din_pass_0_q0 <= cout_drain_IO_L1_out_wrapper372_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper372_U0_fifo_cout_drain_out_V_V_din_pass_0_in = cout_drain_IO_L1_out_wrapper372_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  cout_drain_IO_L1_out_wrapper372_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper372_U0_fifo_cout_drain_out_V_V_write_pass_0_q0 <= cout_drain_IO_L1_out_wrapper372_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper372_U0_fifo_cout_drain_out_V_V_write_pass_0_in = cout_drain_IO_L1_out_wrapper372_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_PE_8_1_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_PE_8_1_V_full_n_pass_0_q0 <= fifo_cout_drain_PE_8_1_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_PE_8_1_V_full_n_pass_0_in = fifo_cout_drain_PE_8_1_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper282_U0_fifo_cin_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper282_U0_fifo_cin_out_V_V_din_pass_0_q0 <= PE_wrapper282_U0_fifo_cin_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper282_U0_fifo_cin_out_V_V_din_pass_0_in = PE_wrapper282_U0_fifo_cin_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper282_U0_fifo_cin_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper282_U0_fifo_cin_out_V_V_write_pass_0_q0 <= PE_wrapper282_U0_fifo_cin_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper282_U0_fifo_cin_out_V_V_write_pass_0_in = PE_wrapper282_U0_fifo_cin_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] w_IO_L2_in146_U0_fifo_w_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    w_IO_L2_in146_U0_fifo_w_out_V_V_din_pass_0_q0 <= w_IO_L2_in146_U0_fifo_w_out_V_V_din_pass_0_out;
  end
  assign w_IO_L2_in146_U0_fifo_w_out_V_V_din_pass_0_in = w_IO_L2_in146_U0_fifo_w_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  w_IO_L2_in146_U0_fifo_w_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    w_IO_L2_in146_U0_fifo_w_out_V_V_write_pass_0_q0 <= w_IO_L2_in146_U0_fifo_w_out_V_V_write_pass_0_out;
  end
  assign w_IO_L2_in146_U0_fifo_w_out_V_V_write_pass_0_in = w_IO_L2_in146_U0_fifo_w_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_PE_12_0_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_PE_12_0_V_full_n_pass_1_q0 <= fifo_cout_drain_PE_12_0_V_full_n_pass_1_out;
  end
  assign fifo_cout_drain_PE_12_0_V_full_n_pass_1_in = fifo_cout_drain_PE_12_0_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_11_1_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_11_1_V_V_full_n_pass_0_q0 <= fifo_cin_PE_11_1_V_V_full_n_pass_0_out;
  end
  assign fifo_cin_PE_11_1_V_V_full_n_pass_0_in = fifo_cin_PE_11_1_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_w_w_IO_L2_in_10_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_w_IO_L2_in_10_V_V_full_n_pass_0_q0 <= fifo_w_w_IO_L2_in_10_V_V_full_n_pass_0_out;
  end
  assign fifo_w_w_IO_L2_in_10_V_V_full_n_pass_0_in = fifo_w_w_IO_L2_in_10_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_cout_drain_IO_L1_out_1_12_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_cout_drain_IO_L1_out_1_12_V_V_full_n_pass_0_q0 <= fifo_cout_drain_cout_drain_IO_L1_out_1_12_V_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_cout_drain_IO_L1_out_1_12_V_V_full_n_pass_0_in = fifo_cout_drain_cout_drain_IO_L1_out_1_12_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg [63:0] cout_drain_IO_L1_out_wrapper404_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper404_U0_fifo_cout_drain_out_V_V_din_pass_0_q0 <= cout_drain_IO_L1_out_wrapper404_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper404_U0_fifo_cout_drain_out_V_V_din_pass_0_in = cout_drain_IO_L1_out_wrapper404_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  cout_drain_IO_L1_out_wrapper404_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper404_U0_fifo_cout_drain_out_V_V_write_pass_0_q0 <= cout_drain_IO_L1_out_wrapper404_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper404_U0_fifo_cout_drain_out_V_V_write_pass_0_in = cout_drain_IO_L1_out_wrapper404_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper283_U0_fifo_cin_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper283_U0_fifo_cin_out_V_V_din_pass_0_q0 <= PE_wrapper283_U0_fifo_cin_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper283_U0_fifo_cin_out_V_V_din_pass_0_in = PE_wrapper283_U0_fifo_cin_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper283_U0_fifo_cin_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper283_U0_fifo_cin_out_V_V_write_pass_0_q0 <= PE_wrapper283_U0_fifo_cin_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper283_U0_fifo_cin_out_V_V_write_pass_0_in = PE_wrapper283_U0_fifo_cin_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_10_0_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_10_0_V_V_full_n_pass_0_q0 <= fifo_cin_PE_10_0_V_V_full_n_pass_0_out;
  end
  assign fifo_cin_PE_10_0_V_V_full_n_pass_0_in = fifo_cin_PE_10_0_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_cout_drain_IO_L1_out_0_13_V_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_cout_drain_IO_L1_out_0_13_V_V_full_n_pass_1_q0 <= fifo_cout_drain_cout_drain_IO_L1_out_0_13_V_V_full_n_pass_1_out;
  end
  assign fifo_cout_drain_cout_drain_IO_L1_out_0_13_V_V_full_n_pass_1_in = fifo_cout_drain_cout_drain_IO_L1_out_0_13_V_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper270_U0_fifo_w_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper270_U0_fifo_w_out_V_V_din_pass_0_q0 <= PE_wrapper270_U0_fifo_w_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper270_U0_fifo_w_out_V_V_din_pass_0_in = PE_wrapper270_U0_fifo_w_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper270_U0_fifo_w_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper270_U0_fifo_w_out_V_V_write_pass_0_q0 <= PE_wrapper270_U0_fifo_w_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper270_U0_fifo_w_out_V_V_write_pass_0_in = PE_wrapper270_U0_fifo_w_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper284_U0_fifo_w_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper284_U0_fifo_w_out_V_V_din_pass_0_q0 <= PE_wrapper284_U0_fifo_w_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper284_U0_fifo_w_out_V_V_din_pass_0_in = PE_wrapper284_U0_fifo_w_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper284_U0_fifo_w_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper284_U0_fifo_w_out_V_V_write_pass_0_q0 <= PE_wrapper284_U0_fifo_w_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper284_U0_fifo_w_out_V_V_write_pass_0_in = PE_wrapper284_U0_fifo_w_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [63:0] cout_drain_IO_L1_out_wrapper390_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper390_U0_fifo_cout_drain_out_V_V_din_pass_0_q0 <= cout_drain_IO_L1_out_wrapper390_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper390_U0_fifo_cout_drain_out_V_V_din_pass_0_in = cout_drain_IO_L1_out_wrapper390_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  cout_drain_IO_L1_out_wrapper390_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper390_U0_fifo_cout_drain_out_V_V_write_pass_0_q0 <= cout_drain_IO_L1_out_wrapper390_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper390_U0_fifo_cout_drain_out_V_V_write_pass_0_in = cout_drain_IO_L1_out_wrapper390_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_PE_9_1_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_PE_9_1_V_full_n_pass_0_q0 <= fifo_cout_drain_PE_9_1_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_PE_9_1_V_full_n_pass_0_in = fifo_cout_drain_PE_9_1_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper272_U0_fifo_w_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper272_U0_fifo_w_out_V_V_din_pass_0_q0 <= PE_wrapper272_U0_fifo_w_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper272_U0_fifo_w_out_V_V_din_pass_0_in = PE_wrapper272_U0_fifo_w_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper272_U0_fifo_w_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper272_U0_fifo_w_out_V_V_write_pass_0_q0 <= PE_wrapper272_U0_fifo_w_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper272_U0_fifo_w_out_V_V_write_pass_0_in = PE_wrapper272_U0_fifo_w_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper284_U0_fifo_cin_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper284_U0_fifo_cin_out_V_V_din_pass_0_q0 <= PE_wrapper284_U0_fifo_cin_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper284_U0_fifo_cin_out_V_V_din_pass_0_in = PE_wrapper284_U0_fifo_cin_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper284_U0_fifo_cin_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper284_U0_fifo_cin_out_V_V_write_pass_0_q0 <= PE_wrapper284_U0_fifo_cin_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper284_U0_fifo_cin_out_V_V_write_pass_0_in = PE_wrapper284_U0_fifo_cin_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_PE_10_1_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_PE_10_1_V_full_n_pass_0_q0 <= fifo_cout_drain_PE_10_1_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_PE_10_1_V_full_n_pass_0_in = fifo_cout_drain_PE_10_1_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  ap_done_Boundary_X0Y2_To_X2Y2_q0;
  always @ (posedge ap_clk) begin
    ap_done_Boundary_X0Y2_To_X2Y2_q0 <= ap_done_Boundary_X0Y2_To_X2Y2_out;
  end
  assign ap_done_Boundary_X0Y2_To_X2Y2_in = ap_done_Boundary_X0Y2_To_X2Y2_q0;
  (* dont_touch = "yes" *) reg  ap_start_Boundary_X0Y4_To_X2Y4_q0;
  always @ (posedge ap_clk) begin
    ap_start_Boundary_X0Y4_To_X2Y4_q0 <= ap_start_Boundary_X0Y4_To_X2Y4_out;
  end
  assign ap_start_Boundary_X0Y4_To_X2Y4_in = ap_start_Boundary_X0Y4_To_X2Y4_q0;
  (* dont_touch = "yes" *) reg  ap_rst_n_Boundary_X0Y4_To_X2Y4_q0;
  always @ (posedge ap_clk) begin
    ap_rst_n_Boundary_X0Y4_To_X2Y4_q0 <= ap_rst_n_Boundary_X0Y4_To_X2Y4_out;
  end
  assign ap_rst_n_Boundary_X0Y4_To_X2Y4_in = ap_rst_n_Boundary_X0Y4_To_X2Y4_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper212_U0_fifo_cin_out_V_V_din_pass_2_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper212_U0_fifo_cin_out_V_V_din_pass_2_q0 <= PE_wrapper212_U0_fifo_cin_out_V_V_din_pass_2_out;
  end
  assign PE_wrapper212_U0_fifo_cin_out_V_V_din_pass_2_in = PE_wrapper212_U0_fifo_cin_out_V_V_din_pass_2_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_6_2_V_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_6_2_V_V_full_n_pass_1_q0 <= fifo_cin_PE_6_2_V_V_full_n_pass_1_out;
  end
  assign fifo_cin_PE_6_2_V_V_full_n_pass_1_in = fifo_cin_PE_6_2_V_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper212_U0_fifo_cin_out_V_V_write_pass_2_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper212_U0_fifo_cin_out_V_V_write_pass_2_q0 <= PE_wrapper212_U0_fifo_cin_out_V_V_write_pass_2_out;
  end
  assign PE_wrapper212_U0_fifo_cin_out_V_V_write_pass_2_in = PE_wrapper212_U0_fifo_cin_out_V_V_write_pass_2_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper213_U0_fifo_cin_out_V_V_din_pass_2_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper213_U0_fifo_cin_out_V_V_din_pass_2_q0 <= PE_wrapper213_U0_fifo_cin_out_V_V_din_pass_2_out;
  end
  assign PE_wrapper213_U0_fifo_cin_out_V_V_din_pass_2_in = PE_wrapper213_U0_fifo_cin_out_V_V_din_pass_2_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_6_3_V_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_6_3_V_V_full_n_pass_1_q0 <= fifo_cin_PE_6_3_V_V_full_n_pass_1_out;
  end
  assign fifo_cin_PE_6_3_V_V_full_n_pass_1_in = fifo_cin_PE_6_3_V_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper213_U0_fifo_cin_out_V_V_write_pass_2_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper213_U0_fifo_cin_out_V_V_write_pass_2_q0 <= PE_wrapper213_U0_fifo_cin_out_V_V_write_pass_2_out;
  end
  assign PE_wrapper213_U0_fifo_cin_out_V_V_write_pass_2_in = PE_wrapper213_U0_fifo_cin_out_V_V_write_pass_2_q0;
  (* dont_touch = "yes" *) reg [63:0] cout_drain_IO_L1_out_wrapper374_U0_fifo_cout_drain_out_V_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper374_U0_fifo_cout_drain_out_V_V_din_pass_1_q0 <= cout_drain_IO_L1_out_wrapper374_U0_fifo_cout_drain_out_V_V_din_pass_1_out;
  end
  assign cout_drain_IO_L1_out_wrapper374_U0_fifo_cout_drain_out_V_V_din_pass_1_in = cout_drain_IO_L1_out_wrapper374_U0_fifo_cout_drain_out_V_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_cout_drain_IO_L1_out_0_8_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_cout_drain_IO_L1_out_0_8_V_V_full_n_pass_0_q0 <= fifo_cout_drain_cout_drain_IO_L1_out_0_8_V_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_cout_drain_IO_L1_out_0_8_V_V_full_n_pass_0_in = fifo_cout_drain_cout_drain_IO_L1_out_0_8_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  cout_drain_IO_L1_out_wrapper374_U0_fifo_cout_drain_out_V_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper374_U0_fifo_cout_drain_out_V_V_write_pass_1_q0 <= cout_drain_IO_L1_out_wrapper374_U0_fifo_cout_drain_out_V_V_write_pass_1_out;
  end
  assign cout_drain_IO_L1_out_wrapper374_U0_fifo_cout_drain_out_V_V_write_pass_1_in = cout_drain_IO_L1_out_wrapper374_U0_fifo_cout_drain_out_V_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_w_w_IO_L2_in_6_V_V_full_n_pass_2_q0;
  always @ (posedge ap_clk) begin
    fifo_w_w_IO_L2_in_6_V_V_full_n_pass_2_q0 <= fifo_w_w_IO_L2_in_6_V_V_full_n_pass_2_out;
  end
  assign fifo_w_w_IO_L2_in_6_V_V_full_n_pass_2_in = fifo_w_w_IO_L2_in_6_V_V_full_n_pass_2_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper260_U0_fifo_cin_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper260_U0_fifo_cin_out_V_V_din_pass_0_q0 <= PE_wrapper260_U0_fifo_cin_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper260_U0_fifo_cin_out_V_V_din_pass_0_in = PE_wrapper260_U0_fifo_cin_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper260_U0_fifo_cin_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper260_U0_fifo_cin_out_V_V_write_pass_0_q0 <= PE_wrapper260_U0_fifo_cin_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper260_U0_fifo_cin_out_V_V_write_pass_0_in = PE_wrapper260_U0_fifo_cin_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_7_2_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_7_2_V_V_full_n_pass_0_q0 <= fifo_cin_PE_7_2_V_V_full_n_pass_0_out;
  end
  assign fifo_cin_PE_7_2_V_V_full_n_pass_0_in = fifo_cin_PE_7_2_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper261_U0_fifo_w_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper261_U0_fifo_w_out_V_V_din_pass_0_q0 <= PE_wrapper261_U0_fifo_w_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper261_U0_fifo_w_out_V_V_din_pass_0_in = PE_wrapper261_U0_fifo_w_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper261_U0_fifo_w_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper261_U0_fifo_w_out_V_V_write_pass_0_q0 <= PE_wrapper261_U0_fifo_w_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper261_U0_fifo_w_out_V_V_write_pass_0_in = PE_wrapper261_U0_fifo_w_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_PE_7_1_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_PE_7_1_V_full_n_pass_0_q0 <= fifo_cout_drain_PE_7_1_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_PE_7_1_V_full_n_pass_0_in = fifo_cout_drain_PE_7_1_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_PE_6_3_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_PE_6_3_V_full_n_pass_0_q0 <= fifo_cout_drain_PE_6_3_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_PE_6_3_V_full_n_pass_0_in = fifo_cout_drain_PE_6_3_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] w_IO_L2_in141_U0_fifo_w_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    w_IO_L2_in141_U0_fifo_w_out_V_V_din_pass_0_q0 <= w_IO_L2_in141_U0_fifo_w_out_V_V_din_pass_0_out;
  end
  assign w_IO_L2_in141_U0_fifo_w_out_V_V_din_pass_0_in = w_IO_L2_in141_U0_fifo_w_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  w_IO_L2_in141_U0_fifo_w_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    w_IO_L2_in141_U0_fifo_w_out_V_V_write_pass_0_q0 <= w_IO_L2_in141_U0_fifo_w_out_V_V_write_pass_0_out;
  end
  assign w_IO_L2_in141_U0_fifo_w_out_V_V_write_pass_0_in = w_IO_L2_in141_U0_fifo_w_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_PE_6_0_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_PE_6_0_V_full_n_pass_0_q0 <= fifo_cout_drain_PE_6_0_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_PE_6_0_V_full_n_pass_0_in = fifo_cout_drain_PE_6_0_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_8_2_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_8_2_V_V_full_n_pass_0_q0 <= fifo_w_PE_8_2_V_V_full_n_pass_0_out;
  end
  assign fifo_w_PE_8_2_V_V_full_n_pass_0_in = fifo_w_PE_8_2_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg [63:0] cout_drain_IO_L1_out_wrapper424_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper424_U0_fifo_cout_drain_out_V_V_din_pass_0_q0 <= cout_drain_IO_L1_out_wrapper424_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper424_U0_fifo_cout_drain_out_V_V_din_pass_0_in = cout_drain_IO_L1_out_wrapper424_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  cout_drain_IO_L1_out_wrapper424_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper424_U0_fifo_cout_drain_out_V_V_write_pass_0_q0 <= cout_drain_IO_L1_out_wrapper424_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper424_U0_fifo_cout_drain_out_V_V_write_pass_0_in = cout_drain_IO_L1_out_wrapper424_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_6_1_V_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_6_1_V_V_full_n_pass_1_q0 <= fifo_cin_PE_6_1_V_V_full_n_pass_1_out;
  end
  assign fifo_cin_PE_6_1_V_V_full_n_pass_1_in = fifo_cin_PE_6_1_V_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_cout_drain_IO_L1_out_3_9_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_cout_drain_IO_L1_out_3_9_V_V_full_n_pass_0_q0 <= fifo_cout_drain_cout_drain_IO_L1_out_3_9_V_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_cout_drain_IO_L1_out_3_9_V_V_full_n_pass_0_in = fifo_cout_drain_cout_drain_IO_L1_out_3_9_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] w_IO_L2_in141_U0_fifo_w_local_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    w_IO_L2_in141_U0_fifo_w_local_out_V_V_din_pass_0_q0 <= w_IO_L2_in141_U0_fifo_w_local_out_V_V_din_pass_0_out;
  end
  assign w_IO_L2_in141_U0_fifo_w_local_out_V_V_din_pass_0_in = w_IO_L2_in141_U0_fifo_w_local_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  w_IO_L2_in141_U0_fifo_w_local_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    w_IO_L2_in141_U0_fifo_w_local_out_V_V_write_pass_0_q0 <= w_IO_L2_in141_U0_fifo_w_local_out_V_V_write_pass_0_out;
  end
  assign w_IO_L2_in141_U0_fifo_w_local_out_V_V_write_pass_0_in = w_IO_L2_in141_U0_fifo_w_local_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [31:0] PE_wrapper261_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper261_U0_fifo_cout_drain_out_V_din_pass_0_q0 <= PE_wrapper261_U0_fifo_cout_drain_out_V_din_pass_0_out;
  end
  assign PE_wrapper261_U0_fifo_cout_drain_out_V_din_pass_0_in = PE_wrapper261_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper261_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper261_U0_fifo_cout_drain_out_V_write_pass_0_q0 <= PE_wrapper261_U0_fifo_cout_drain_out_V_write_pass_0_out;
  end
  assign PE_wrapper261_U0_fifo_cout_drain_out_V_write_pass_0_in = PE_wrapper261_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_6_1_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_6_1_V_V_full_n_pass_0_q0 <= fifo_w_PE_6_1_V_V_full_n_pass_0_out;
  end
  assign fifo_w_PE_6_1_V_V_full_n_pass_0_in = fifo_w_PE_6_1_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg [63:0] cout_drain_IO_L1_out_wrapper376_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper376_U0_fifo_cout_drain_out_V_V_din_pass_0_q0 <= cout_drain_IO_L1_out_wrapper376_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper376_U0_fifo_cout_drain_out_V_V_din_pass_0_in = cout_drain_IO_L1_out_wrapper376_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  cout_drain_IO_L1_out_wrapper376_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper376_U0_fifo_cout_drain_out_V_V_write_pass_0_q0 <= cout_drain_IO_L1_out_wrapper376_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper376_U0_fifo_cout_drain_out_V_V_write_pass_0_in = cout_drain_IO_L1_out_wrapper376_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper236_U0_fifo_w_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper236_U0_fifo_w_out_V_V_din_pass_0_q0 <= PE_wrapper236_U0_fifo_w_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper236_U0_fifo_w_out_V_V_din_pass_0_in = PE_wrapper236_U0_fifo_w_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper236_U0_fifo_w_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper236_U0_fifo_w_out_V_V_write_pass_0_q0 <= PE_wrapper236_U0_fifo_w_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper236_U0_fifo_w_out_V_V_write_pass_0_in = PE_wrapper236_U0_fifo_w_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper223_U0_fifo_cin_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper223_U0_fifo_cin_out_V_V_din_pass_0_q0 <= PE_wrapper223_U0_fifo_cin_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper223_U0_fifo_cin_out_V_V_din_pass_0_in = PE_wrapper223_U0_fifo_cin_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper223_U0_fifo_cin_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper223_U0_fifo_cin_out_V_V_write_pass_0_q0 <= PE_wrapper223_U0_fifo_cin_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper223_U0_fifo_cin_out_V_V_write_pass_0_in = PE_wrapper223_U0_fifo_cin_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_cout_drain_IO_L1_out_2_10_V_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_cout_drain_IO_L1_out_2_10_V_V_full_n_pass_1_q0 <= fifo_cout_drain_cout_drain_IO_L1_out_2_10_V_V_full_n_pass_1_out;
  end
  assign fifo_cout_drain_cout_drain_IO_L1_out_2_10_V_V_full_n_pass_1_in = fifo_cout_drain_cout_drain_IO_L1_out_2_10_V_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper249_U0_fifo_w_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper249_U0_fifo_w_out_V_V_din_pass_0_q0 <= PE_wrapper249_U0_fifo_w_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper249_U0_fifo_w_out_V_V_din_pass_0_in = PE_wrapper249_U0_fifo_w_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper249_U0_fifo_w_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper249_U0_fifo_w_out_V_V_write_pass_0_q0 <= PE_wrapper249_U0_fifo_w_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper249_U0_fifo_w_out_V_V_write_pass_0_in = PE_wrapper249_U0_fifo_w_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper223_U0_fifo_w_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper223_U0_fifo_w_out_V_V_din_pass_0_q0 <= PE_wrapper223_U0_fifo_w_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper223_U0_fifo_w_out_V_V_din_pass_0_in = PE_wrapper223_U0_fifo_w_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper223_U0_fifo_w_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper223_U0_fifo_w_out_V_V_write_pass_0_q0 <= PE_wrapper223_U0_fifo_w_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper223_U0_fifo_w_out_V_V_write_pass_0_in = PE_wrapper223_U0_fifo_w_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_9_2_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_9_2_V_V_full_n_pass_0_q0 <= fifo_w_PE_9_2_V_V_full_n_pass_0_out;
  end
  assign fifo_w_PE_9_2_V_V_full_n_pass_0_in = fifo_w_PE_9_2_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_cout_drain_IO_L1_out_1_8_V_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_cout_drain_IO_L1_out_1_8_V_V_full_n_pass_1_q0 <= fifo_cout_drain_cout_drain_IO_L1_out_1_8_V_V_full_n_pass_1_out;
  end
  assign fifo_cout_drain_cout_drain_IO_L1_out_1_8_V_V_full_n_pass_1_in = fifo_cout_drain_cout_drain_IO_L1_out_1_8_V_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_8_3_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_8_3_V_V_full_n_pass_0_q0 <= fifo_cin_PE_8_3_V_V_full_n_pass_0_out;
  end
  assign fifo_cin_PE_8_3_V_V_full_n_pass_0_in = fifo_cin_PE_8_3_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg [63:0] cout_drain_IO_L1_out_wrapper408_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper408_U0_fifo_cout_drain_out_V_V_din_pass_0_q0 <= cout_drain_IO_L1_out_wrapper408_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper408_U0_fifo_cout_drain_out_V_V_din_pass_0_in = cout_drain_IO_L1_out_wrapper408_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  cout_drain_IO_L1_out_wrapper408_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper408_U0_fifo_cout_drain_out_V_V_write_pass_0_q0 <= cout_drain_IO_L1_out_wrapper408_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper408_U0_fifo_cout_drain_out_V_V_write_pass_0_in = cout_drain_IO_L1_out_wrapper408_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_PE_6_2_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_PE_6_2_V_full_n_pass_0_q0 <= fifo_cout_drain_PE_6_2_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_PE_6_2_V_full_n_pass_0_in = fifo_cout_drain_PE_6_2_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_7_2_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_7_2_V_V_full_n_pass_0_q0 <= fifo_w_PE_7_2_V_V_full_n_pass_0_out;
  end
  assign fifo_w_PE_7_2_V_V_full_n_pass_0_in = fifo_w_PE_7_2_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper261_U0_fifo_cin_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper261_U0_fifo_cin_out_V_V_din_pass_0_q0 <= PE_wrapper261_U0_fifo_cin_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper261_U0_fifo_cin_out_V_V_din_pass_0_in = PE_wrapper261_U0_fifo_cin_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper261_U0_fifo_cin_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper261_U0_fifo_cin_out_V_V_write_pass_0_q0 <= PE_wrapper261_U0_fifo_cin_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper261_U0_fifo_cin_out_V_V_write_pass_0_in = PE_wrapper261_U0_fifo_cin_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_cout_drain_IO_L1_out_0_7_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_cout_drain_IO_L1_out_0_7_V_V_full_n_pass_0_q0 <= fifo_cout_drain_cout_drain_IO_L1_out_0_7_V_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_cout_drain_IO_L1_out_0_7_V_V_full_n_pass_0_in = fifo_cout_drain_cout_drain_IO_L1_out_0_7_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg [63:0] cout_drain_IO_L1_out_wrapper392_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper392_U0_fifo_cout_drain_out_V_V_din_pass_0_q0 <= cout_drain_IO_L1_out_wrapper392_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper392_U0_fifo_cout_drain_out_V_V_din_pass_0_in = cout_drain_IO_L1_out_wrapper392_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  cout_drain_IO_L1_out_wrapper392_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper392_U0_fifo_cout_drain_out_V_V_write_pass_0_q0 <= cout_drain_IO_L1_out_wrapper392_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper392_U0_fifo_cout_drain_out_V_V_write_pass_0_in = cout_drain_IO_L1_out_wrapper392_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_PE_7_3_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_PE_7_3_V_full_n_pass_0_q0 <= fifo_cout_drain_PE_7_3_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_PE_7_3_V_full_n_pass_0_in = fifo_cout_drain_PE_7_3_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  ap_done_Boundary_X4Y0_To_X4Y2_q0;
  always @ (posedge ap_clk) begin
    ap_done_Boundary_X4Y0_To_X4Y2_q0 <= ap_done_Boundary_X4Y0_To_X4Y2_out;
  end
  assign ap_done_Boundary_X4Y0_To_X4Y2_in = ap_done_Boundary_X4Y0_To_X4Y2_q0;
  (* dont_touch = "yes" *) reg  ap_start_Boundary_X2Y2_To_X4Y2_q0;
  always @ (posedge ap_clk) begin
    ap_start_Boundary_X2Y2_To_X4Y2_q0 <= ap_start_Boundary_X2Y2_To_X4Y2_out;
  end
  assign ap_start_Boundary_X2Y2_To_X4Y2_in = ap_start_Boundary_X2Y2_To_X4Y2_q0;
  (* dont_touch = "yes" *) reg  ap_rst_n_Boundary_X2Y2_To_X4Y2_q0;
  always @ (posedge ap_clk) begin
    ap_rst_n_Boundary_X2Y2_To_X4Y2_q0 <= ap_rst_n_Boundary_X2Y2_To_X4Y2_out;
  end
  assign ap_rst_n_Boundary_X2Y2_To_X4Y2_in = ap_rst_n_Boundary_X2Y2_To_X4Y2_q0;
  (* dont_touch = "yes" *) reg  ap_start_Boundary_X2Y0_To_X2Y2_q0;
  always @ (posedge ap_clk) begin
    ap_start_Boundary_X2Y0_To_X2Y2_q0 <= ap_start_Boundary_X2Y0_To_X2Y2_out;
  end
  assign ap_start_Boundary_X2Y0_To_X2Y2_in = ap_start_Boundary_X2Y0_To_X2Y2_q0;
  (* dont_touch = "yes" *) reg  ap_rst_n_Boundary_X2Y0_To_X2Y2_q0;
  always @ (posedge ap_clk) begin
    ap_rst_n_Boundary_X2Y0_To_X2Y2_q0 <= ap_rst_n_Boundary_X2Y0_To_X2Y2_out;
  end
  assign ap_rst_n_Boundary_X2Y0_To_X2Y2_in = ap_rst_n_Boundary_X2Y0_To_X2Y2_q0;
  (* dont_touch = "yes" *) reg [255:0] w_IO_L2_in140_U0_fifo_w_out_V_V_din_pass_2_q0;
  always @ (posedge ap_clk) begin
    w_IO_L2_in140_U0_fifo_w_out_V_V_din_pass_2_q0 <= w_IO_L2_in140_U0_fifo_w_out_V_V_din_pass_2_out;
  end
  assign w_IO_L2_in140_U0_fifo_w_out_V_V_din_pass_2_in = w_IO_L2_in140_U0_fifo_w_out_V_V_din_pass_2_q0;
  (* dont_touch = "yes" *) reg  fifo_w_w_IO_L2_in_6_V_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_w_w_IO_L2_in_6_V_V_full_n_pass_1_q0 <= fifo_w_w_IO_L2_in_6_V_V_full_n_pass_1_out;
  end
  assign fifo_w_w_IO_L2_in_6_V_V_full_n_pass_1_in = fifo_w_w_IO_L2_in_6_V_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg  w_IO_L2_in140_U0_fifo_w_out_V_V_write_pass_2_q0;
  always @ (posedge ap_clk) begin
    w_IO_L2_in140_U0_fifo_w_out_V_V_write_pass_2_q0 <= w_IO_L2_in140_U0_fifo_w_out_V_V_write_pass_2_out;
  end
  assign w_IO_L2_in140_U0_fifo_w_out_V_V_write_pass_2_in = w_IO_L2_in140_U0_fifo_w_out_V_V_write_pass_2_q0;
  (* dont_touch = "yes" *) reg [63:0] cout_drain_IO_L1_out_wrapper404_U0_fifo_cout_drain_out_V_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper404_U0_fifo_cout_drain_out_V_V_din_pass_1_q0 <= cout_drain_IO_L1_out_wrapper404_U0_fifo_cout_drain_out_V_V_din_pass_1_out;
  end
  assign cout_drain_IO_L1_out_wrapper404_U0_fifo_cout_drain_out_V_V_din_pass_1_in = cout_drain_IO_L1_out_wrapper404_U0_fifo_cout_drain_out_V_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_cout_drain_IO_L1_out_2_10_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_cout_drain_IO_L1_out_2_10_V_V_full_n_pass_0_q0 <= fifo_cout_drain_cout_drain_IO_L1_out_2_10_V_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_cout_drain_IO_L1_out_2_10_V_V_full_n_pass_0_in = fifo_cout_drain_cout_drain_IO_L1_out_2_10_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  cout_drain_IO_L1_out_wrapper404_U0_fifo_cout_drain_out_V_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper404_U0_fifo_cout_drain_out_V_V_write_pass_1_q0 <= cout_drain_IO_L1_out_wrapper404_U0_fifo_cout_drain_out_V_V_write_pass_1_out;
  end
  assign cout_drain_IO_L1_out_wrapper404_U0_fifo_cout_drain_out_V_V_write_pass_1_in = cout_drain_IO_L1_out_wrapper404_U0_fifo_cout_drain_out_V_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [63:0] cout_drain_IO_L1_out_wrapper390_U0_fifo_cout_drain_out_V_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper390_U0_fifo_cout_drain_out_V_V_din_pass_1_q0 <= cout_drain_IO_L1_out_wrapper390_U0_fifo_cout_drain_out_V_V_din_pass_1_out;
  end
  assign cout_drain_IO_L1_out_wrapper390_U0_fifo_cout_drain_out_V_V_din_pass_1_in = cout_drain_IO_L1_out_wrapper390_U0_fifo_cout_drain_out_V_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_cout_drain_IO_L1_out_1_8_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_cout_drain_IO_L1_out_1_8_V_V_full_n_pass_0_q0 <= fifo_cout_drain_cout_drain_IO_L1_out_1_8_V_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_cout_drain_IO_L1_out_1_8_V_V_full_n_pass_0_in = fifo_cout_drain_cout_drain_IO_L1_out_1_8_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  cout_drain_IO_L1_out_wrapper390_U0_fifo_cout_drain_out_V_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper390_U0_fifo_cout_drain_out_V_V_write_pass_1_q0 <= cout_drain_IO_L1_out_wrapper390_U0_fifo_cout_drain_out_V_V_write_pass_1_out;
  end
  assign cout_drain_IO_L1_out_wrapper390_U0_fifo_cout_drain_out_V_V_write_pass_1_in = cout_drain_IO_L1_out_wrapper390_U0_fifo_cout_drain_out_V_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper249_U0_fifo_w_out_V_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper249_U0_fifo_w_out_V_V_din_pass_1_q0 <= PE_wrapper249_U0_fifo_w_out_V_V_din_pass_1_out;
  end
  assign PE_wrapper249_U0_fifo_w_out_V_V_din_pass_1_in = PE_wrapper249_U0_fifo_w_out_V_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_8_4_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_8_4_V_V_full_n_pass_0_q0 <= fifo_w_PE_8_4_V_V_full_n_pass_0_out;
  end
  assign fifo_w_PE_8_4_V_V_full_n_pass_0_in = fifo_w_PE_8_4_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper249_U0_fifo_w_out_V_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper249_U0_fifo_w_out_V_V_write_pass_1_q0 <= PE_wrapper249_U0_fifo_w_out_V_V_write_pass_1_out;
  end
  assign PE_wrapper249_U0_fifo_w_out_V_V_write_pass_1_in = PE_wrapper249_U0_fifo_w_out_V_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper272_U0_fifo_w_out_V_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper272_U0_fifo_w_out_V_V_din_pass_1_q0 <= PE_wrapper272_U0_fifo_w_out_V_V_din_pass_1_out;
  end
  assign PE_wrapper272_U0_fifo_w_out_V_V_din_pass_1_in = PE_wrapper272_U0_fifo_w_out_V_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_10_3_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_10_3_V_V_full_n_pass_0_q0 <= fifo_w_PE_10_3_V_V_full_n_pass_0_out;
  end
  assign fifo_w_PE_10_3_V_V_full_n_pass_0_in = fifo_w_PE_10_3_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper272_U0_fifo_w_out_V_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper272_U0_fifo_w_out_V_V_write_pass_1_q0 <= PE_wrapper272_U0_fifo_w_out_V_V_write_pass_1_out;
  end
  assign PE_wrapper272_U0_fifo_w_out_V_V_write_pass_1_in = PE_wrapper272_U0_fifo_w_out_V_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper261_U0_fifo_cin_out_V_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper261_U0_fifo_cin_out_V_V_din_pass_1_q0 <= PE_wrapper261_U0_fifo_cin_out_V_V_din_pass_1_out;
  end
  assign PE_wrapper261_U0_fifo_cin_out_V_V_din_pass_1_in = PE_wrapper261_U0_fifo_cin_out_V_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_10_3_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_10_3_V_V_full_n_pass_0_q0 <= fifo_cin_PE_10_3_V_V_full_n_pass_0_out;
  end
  assign fifo_cin_PE_10_3_V_V_full_n_pass_0_in = fifo_cin_PE_10_3_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper261_U0_fifo_cin_out_V_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper261_U0_fifo_cin_out_V_V_write_pass_1_q0 <= PE_wrapper261_U0_fifo_cin_out_V_V_write_pass_1_out;
  end
  assign PE_wrapper261_U0_fifo_cin_out_V_V_write_pass_1_in = PE_wrapper261_U0_fifo_cin_out_V_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper224_U0_fifo_cin_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper224_U0_fifo_cin_out_V_V_din_pass_0_q0 <= PE_wrapper224_U0_fifo_cin_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper224_U0_fifo_cin_out_V_V_din_pass_0_in = PE_wrapper224_U0_fifo_cin_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper224_U0_fifo_cin_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper224_U0_fifo_cin_out_V_V_write_pass_0_q0 <= PE_wrapper224_U0_fifo_cin_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper224_U0_fifo_cin_out_V_V_write_pass_0_in = PE_wrapper224_U0_fifo_cin_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [31:0] PE_wrapper235_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper235_U0_fifo_cout_drain_out_V_din_pass_0_q0 <= PE_wrapper235_U0_fifo_cout_drain_out_V_din_pass_0_out;
  end
  assign PE_wrapper235_U0_fifo_cout_drain_out_V_din_pass_0_in = PE_wrapper235_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper235_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper235_U0_fifo_cout_drain_out_V_write_pass_0_q0 <= PE_wrapper235_U0_fifo_cout_drain_out_V_write_pass_0_out;
  end
  assign PE_wrapper235_U0_fifo_cout_drain_out_V_write_pass_0_in = PE_wrapper235_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [31:0] PE_wrapper225_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper225_U0_fifo_cout_drain_out_V_din_pass_0_q0 <= PE_wrapper225_U0_fifo_cout_drain_out_V_din_pass_0_out;
  end
  assign PE_wrapper225_U0_fifo_cout_drain_out_V_din_pass_0_in = PE_wrapper225_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper225_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper225_U0_fifo_cout_drain_out_V_write_pass_0_q0 <= PE_wrapper225_U0_fifo_cout_drain_out_V_write_pass_0_out;
  end
  assign PE_wrapper225_U0_fifo_cout_drain_out_V_write_pass_0_in = PE_wrapper225_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_w_w_IO_L2_in_7_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_w_IO_L2_in_7_V_V_full_n_pass_0_q0 <= fifo_w_w_IO_L2_in_7_V_V_full_n_pass_0_out;
  end
  assign fifo_w_w_IO_L2_in_7_V_V_full_n_pass_0_in = fifo_w_w_IO_L2_in_7_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper235_U0_fifo_cin_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper235_U0_fifo_cin_out_V_V_din_pass_0_q0 <= PE_wrapper235_U0_fifo_cin_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper235_U0_fifo_cin_out_V_V_din_pass_0_in = PE_wrapper235_U0_fifo_cin_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper235_U0_fifo_cin_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper235_U0_fifo_cin_out_V_V_write_pass_0_q0 <= PE_wrapper235_U0_fifo_cin_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper235_U0_fifo_cin_out_V_V_write_pass_0_in = PE_wrapper235_U0_fifo_cin_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [31:0] PE_wrapper222_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper222_U0_fifo_cout_drain_out_V_din_pass_0_q0 <= PE_wrapper222_U0_fifo_cout_drain_out_V_din_pass_0_out;
  end
  assign PE_wrapper222_U0_fifo_cout_drain_out_V_din_pass_0_in = PE_wrapper222_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper222_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper222_U0_fifo_cout_drain_out_V_write_pass_0_q0 <= PE_wrapper222_U0_fifo_cout_drain_out_V_write_pass_0_out;
  end
  assign PE_wrapper222_U0_fifo_cout_drain_out_V_write_pass_0_in = PE_wrapper222_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_6_2_V_V_full_n_pass_2_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_6_2_V_V_full_n_pass_2_q0 <= fifo_cin_PE_6_2_V_V_full_n_pass_2_out;
  end
  assign fifo_cin_PE_6_2_V_V_full_n_pass_2_in = fifo_cin_PE_6_2_V_V_full_n_pass_2_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper225_U0_fifo_w_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper225_U0_fifo_w_out_V_V_din_pass_0_q0 <= PE_wrapper225_U0_fifo_w_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper225_U0_fifo_w_out_V_V_din_pass_0_in = PE_wrapper225_U0_fifo_w_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper225_U0_fifo_w_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper225_U0_fifo_w_out_V_V_write_pass_0_q0 <= PE_wrapper225_U0_fifo_w_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper225_U0_fifo_w_out_V_V_write_pass_0_in = PE_wrapper225_U0_fifo_w_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [63:0] cout_drain_IO_L1_out_wrapper421_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper421_U0_fifo_cout_drain_out_V_V_din_pass_0_q0 <= cout_drain_IO_L1_out_wrapper421_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper421_U0_fifo_cout_drain_out_V_V_din_pass_0_in = cout_drain_IO_L1_out_wrapper421_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  cout_drain_IO_L1_out_wrapper421_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper421_U0_fifo_cout_drain_out_V_V_write_pass_0_q0 <= cout_drain_IO_L1_out_wrapper421_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper421_U0_fifo_cout_drain_out_V_V_write_pass_0_in = cout_drain_IO_L1_out_wrapper421_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_6_0_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_6_0_V_V_full_n_pass_0_q0 <= fifo_w_PE_6_0_V_V_full_n_pass_0_out;
  end
  assign fifo_w_PE_6_0_V_V_full_n_pass_0_in = fifo_w_PE_6_0_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg [63:0] cout_drain_IO_L1_out_wrapper375_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper375_U0_fifo_cout_drain_out_V_V_din_pass_0_q0 <= cout_drain_IO_L1_out_wrapper375_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper375_U0_fifo_cout_drain_out_V_V_din_pass_0_in = cout_drain_IO_L1_out_wrapper375_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  cout_drain_IO_L1_out_wrapper375_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper375_U0_fifo_cout_drain_out_V_V_write_pass_0_q0 <= cout_drain_IO_L1_out_wrapper375_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper375_U0_fifo_cout_drain_out_V_V_write_pass_0_in = cout_drain_IO_L1_out_wrapper375_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_PE_9_3_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_PE_9_3_V_full_n_pass_0_q0 <= fifo_cout_drain_PE_9_3_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_PE_9_3_V_full_n_pass_0_in = fifo_cout_drain_PE_9_3_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_6_3_V_V_full_n_pass_2_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_6_3_V_V_full_n_pass_2_q0 <= fifo_cin_PE_6_3_V_V_full_n_pass_2_out;
  end
  assign fifo_cin_PE_6_3_V_V_full_n_pass_2_in = fifo_cin_PE_6_3_V_V_full_n_pass_2_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper222_U0_fifo_w_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper222_U0_fifo_w_out_V_V_din_pass_0_q0 <= PE_wrapper222_U0_fifo_w_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper222_U0_fifo_w_out_V_V_din_pass_0_in = PE_wrapper222_U0_fifo_w_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper222_U0_fifo_w_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper222_U0_fifo_w_out_V_V_write_pass_0_q0 <= PE_wrapper222_U0_fifo_w_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper222_U0_fifo_w_out_V_V_write_pass_0_in = PE_wrapper222_U0_fifo_w_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper237_U0_fifo_w_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper237_U0_fifo_w_out_V_V_din_pass_0_q0 <= PE_wrapper237_U0_fifo_w_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper237_U0_fifo_w_out_V_V_din_pass_0_in = PE_wrapper237_U0_fifo_w_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper237_U0_fifo_w_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper237_U0_fifo_w_out_V_V_write_pass_0_q0 <= PE_wrapper237_U0_fifo_w_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper237_U0_fifo_w_out_V_V_write_pass_0_in = PE_wrapper237_U0_fifo_w_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_7_3_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_7_3_V_V_full_n_pass_0_q0 <= fifo_w_PE_7_3_V_V_full_n_pass_0_out;
  end
  assign fifo_w_PE_7_3_V_V_full_n_pass_0_in = fifo_w_PE_7_3_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_7_1_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_7_1_V_V_full_n_pass_0_q0 <= fifo_cin_PE_7_1_V_V_full_n_pass_0_out;
  end
  assign fifo_cin_PE_7_1_V_V_full_n_pass_0_in = fifo_cin_PE_7_1_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_cout_drain_IO_L1_out_0_8_V_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_cout_drain_IO_L1_out_0_8_V_V_full_n_pass_1_q0 <= fifo_cout_drain_cout_drain_IO_L1_out_0_8_V_V_full_n_pass_1_out;
  end
  assign fifo_cout_drain_cout_drain_IO_L1_out_0_8_V_V_full_n_pass_1_in = fifo_cout_drain_cout_drain_IO_L1_out_0_8_V_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_6_2_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_6_2_V_V_full_n_pass_0_q0 <= fifo_w_PE_6_2_V_V_full_n_pass_0_out;
  end
  assign fifo_w_PE_6_2_V_V_full_n_pass_0_in = fifo_w_PE_6_2_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_cout_drain_IO_L1_out_3_10_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_cout_drain_IO_L1_out_3_10_V_V_full_n_pass_0_q0 <= fifo_cout_drain_cout_drain_IO_L1_out_3_10_V_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_cout_drain_IO_L1_out_3_10_V_V_full_n_pass_0_in = fifo_cout_drain_cout_drain_IO_L1_out_3_10_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper234_U0_fifo_cin_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper234_U0_fifo_cin_out_V_V_din_pass_0_q0 <= PE_wrapper234_U0_fifo_cin_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper234_U0_fifo_cin_out_V_V_din_pass_0_in = PE_wrapper234_U0_fifo_cin_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper234_U0_fifo_cin_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper234_U0_fifo_cin_out_V_V_write_pass_0_q0 <= PE_wrapper234_U0_fifo_cin_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper234_U0_fifo_cin_out_V_V_write_pass_0_in = PE_wrapper234_U0_fifo_cin_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper237_U0_fifo_cin_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper237_U0_fifo_cin_out_V_V_din_pass_0_q0 <= PE_wrapper237_U0_fifo_cin_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper237_U0_fifo_cin_out_V_V_din_pass_0_in = PE_wrapper237_U0_fifo_cin_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper237_U0_fifo_cin_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper237_U0_fifo_cin_out_V_V_write_pass_0_q0 <= PE_wrapper237_U0_fifo_cin_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper237_U0_fifo_cin_out_V_V_write_pass_0_in = PE_wrapper237_U0_fifo_cin_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper235_U0_fifo_w_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper235_U0_fifo_w_out_V_V_din_pass_0_q0 <= PE_wrapper235_U0_fifo_w_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper235_U0_fifo_w_out_V_V_din_pass_0_in = PE_wrapper235_U0_fifo_w_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper235_U0_fifo_w_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper235_U0_fifo_w_out_V_V_write_pass_0_q0 <= PE_wrapper235_U0_fifo_w_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper235_U0_fifo_w_out_V_V_write_pass_0_in = PE_wrapper235_U0_fifo_w_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] w_IO_L2_in142_U0_fifo_w_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    w_IO_L2_in142_U0_fifo_w_out_V_V_din_pass_0_q0 <= w_IO_L2_in142_U0_fifo_w_out_V_V_din_pass_0_out;
  end
  assign w_IO_L2_in142_U0_fifo_w_out_V_V_din_pass_0_in = w_IO_L2_in142_U0_fifo_w_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  w_IO_L2_in142_U0_fifo_w_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    w_IO_L2_in142_U0_fifo_w_out_V_V_write_pass_0_q0 <= w_IO_L2_in142_U0_fifo_w_out_V_V_write_pass_0_out;
  end
  assign w_IO_L2_in142_U0_fifo_w_out_V_V_write_pass_0_in = w_IO_L2_in142_U0_fifo_w_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [31:0] PE_wrapper224_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper224_U0_fifo_cout_drain_out_V_din_pass_0_q0 <= PE_wrapper224_U0_fifo_cout_drain_out_V_din_pass_0_out;
  end
  assign PE_wrapper224_U0_fifo_cout_drain_out_V_din_pass_0_in = PE_wrapper224_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper224_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper224_U0_fifo_cout_drain_out_V_write_pass_0_q0 <= PE_wrapper224_U0_fifo_cout_drain_out_V_write_pass_0_out;
  end
  assign PE_wrapper224_U0_fifo_cout_drain_out_V_write_pass_0_in = PE_wrapper224_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_6_0_V_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_6_0_V_V_full_n_pass_1_q0 <= fifo_cin_PE_6_0_V_V_full_n_pass_1_out;
  end
  assign fifo_cin_PE_6_0_V_V_full_n_pass_1_in = fifo_cin_PE_6_0_V_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg [31:0] PE_wrapper237_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper237_U0_fifo_cout_drain_out_V_din_pass_0_q0 <= PE_wrapper237_U0_fifo_cout_drain_out_V_din_pass_0_out;
  end
  assign PE_wrapper237_U0_fifo_cout_drain_out_V_din_pass_0_in = PE_wrapper237_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper237_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper237_U0_fifo_cout_drain_out_V_write_pass_0_q0 <= PE_wrapper237_U0_fifo_cout_drain_out_V_write_pass_0_out;
  end
  assign PE_wrapper237_U0_fifo_cout_drain_out_V_write_pass_0_in = PE_wrapper237_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  ap_done_Boundary_X2Y2_To_X4Y2_q0;
  always @ (posedge ap_clk) begin
    ap_done_Boundary_X2Y2_To_X4Y2_q0 <= ap_done_Boundary_X2Y2_To_X4Y2_out;
  end
  assign ap_done_Boundary_X2Y2_To_X4Y2_in = ap_done_Boundary_X2Y2_To_X4Y2_q0;
  (* dont_touch = "yes" *) reg  ap_start_Boundary_X2Y4_To_X4Y4_q0;
  always @ (posedge ap_clk) begin
    ap_start_Boundary_X2Y4_To_X4Y4_q0 <= ap_start_Boundary_X2Y4_To_X4Y4_out;
  end
  assign ap_start_Boundary_X2Y4_To_X4Y4_in = ap_start_Boundary_X2Y4_To_X4Y4_q0;
  (* dont_touch = "yes" *) reg  ap_rst_n_Boundary_X2Y4_To_X4Y4_q0;
  always @ (posedge ap_clk) begin
    ap_rst_n_Boundary_X2Y4_To_X4Y4_q0 <= ap_rst_n_Boundary_X2Y4_To_X4Y4_out;
  end
  assign ap_rst_n_Boundary_X2Y4_To_X4Y4_in = ap_rst_n_Boundary_X2Y4_To_X4Y4_q0;
  (* dont_touch = "yes" *) reg [63:0] cout_drain_IO_L1_out_wrapper402_U0_fifo_cout_drain_out_V_V_din_pass_2_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper402_U0_fifo_cout_drain_out_V_V_din_pass_2_q0 <= cout_drain_IO_L1_out_wrapper402_U0_fifo_cout_drain_out_V_V_din_pass_2_out;
  end
  assign cout_drain_IO_L1_out_wrapper402_U0_fifo_cout_drain_out_V_V_din_pass_2_in = cout_drain_IO_L1_out_wrapper402_U0_fifo_cout_drain_out_V_V_din_pass_2_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_cout_drain_IO_L1_out_2_12_V_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_cout_drain_IO_L1_out_2_12_V_V_full_n_pass_1_q0 <= fifo_cout_drain_cout_drain_IO_L1_out_2_12_V_V_full_n_pass_1_out;
  end
  assign fifo_cout_drain_cout_drain_IO_L1_out_2_12_V_V_full_n_pass_1_in = fifo_cout_drain_cout_drain_IO_L1_out_2_12_V_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg  cout_drain_IO_L1_out_wrapper402_U0_fifo_cout_drain_out_V_V_write_pass_2_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper402_U0_fifo_cout_drain_out_V_V_write_pass_2_q0 <= cout_drain_IO_L1_out_wrapper402_U0_fifo_cout_drain_out_V_V_write_pass_2_out;
  end
  assign cout_drain_IO_L1_out_wrapper402_U0_fifo_cout_drain_out_V_V_write_pass_2_in = cout_drain_IO_L1_out_wrapper402_U0_fifo_cout_drain_out_V_V_write_pass_2_q0;
  (* dont_touch = "yes" *) reg [31:0] PE_wrapper294_U0_fifo_cout_drain_out_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper294_U0_fifo_cout_drain_out_V_din_pass_1_q0 <= PE_wrapper294_U0_fifo_cout_drain_out_V_din_pass_1_out;
  end
  assign PE_wrapper294_U0_fifo_cout_drain_out_V_din_pass_1_in = PE_wrapper294_U0_fifo_cout_drain_out_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_PE_12_0_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_PE_12_0_V_full_n_pass_0_q0 <= fifo_cout_drain_PE_12_0_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_PE_12_0_V_full_n_pass_0_in = fifo_cout_drain_PE_12_0_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper294_U0_fifo_cout_drain_out_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper294_U0_fifo_cout_drain_out_V_write_pass_1_q0 <= PE_wrapper294_U0_fifo_cout_drain_out_V_write_pass_1_out;
  end
  assign PE_wrapper294_U0_fifo_cout_drain_out_V_write_pass_1_in = PE_wrapper294_U0_fifo_cout_drain_out_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [63:0] cout_drain_IO_L1_out_wrapper369_U0_fifo_cout_drain_out_V_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper369_U0_fifo_cout_drain_out_V_V_din_pass_1_q0 <= cout_drain_IO_L1_out_wrapper369_U0_fifo_cout_drain_out_V_V_din_pass_1_out;
  end
  assign cout_drain_IO_L1_out_wrapper369_U0_fifo_cout_drain_out_V_V_din_pass_1_in = cout_drain_IO_L1_out_wrapper369_U0_fifo_cout_drain_out_V_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_cout_drain_IO_L1_out_0_13_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_cout_drain_IO_L1_out_0_13_V_V_full_n_pass_0_q0 <= fifo_cout_drain_cout_drain_IO_L1_out_0_13_V_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_cout_drain_IO_L1_out_0_13_V_V_full_n_pass_0_in = fifo_cout_drain_cout_drain_IO_L1_out_0_13_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  cout_drain_IO_L1_out_wrapper369_U0_fifo_cout_drain_out_V_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper369_U0_fifo_cout_drain_out_V_V_write_pass_1_q0 <= cout_drain_IO_L1_out_wrapper369_U0_fifo_cout_drain_out_V_V_write_pass_1_out;
  end
  assign cout_drain_IO_L1_out_wrapper369_U0_fifo_cout_drain_out_V_V_write_pass_1_in = cout_drain_IO_L1_out_wrapper369_U0_fifo_cout_drain_out_V_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper298_U0_fifo_cin_out_V_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper298_U0_fifo_cin_out_V_V_din_pass_1_q0 <= PE_wrapper298_U0_fifo_cin_out_V_V_din_pass_1_out;
  end
  assign PE_wrapper298_U0_fifo_cin_out_V_V_din_pass_1_in = PE_wrapper298_U0_fifo_cin_out_V_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_13_4_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_13_4_V_V_full_n_pass_0_q0 <= fifo_cin_PE_13_4_V_V_full_n_pass_0_out;
  end
  assign fifo_cin_PE_13_4_V_V_full_n_pass_0_in = fifo_cin_PE_13_4_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper298_U0_fifo_cin_out_V_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper298_U0_fifo_cin_out_V_V_write_pass_1_q0 <= PE_wrapper298_U0_fifo_cin_out_V_V_write_pass_1_out;
  end
  assign PE_wrapper298_U0_fifo_cin_out_V_V_write_pass_1_in = PE_wrapper298_U0_fifo_cin_out_V_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [31:0] PE_wrapper250_U0_fifo_cout_drain_out_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper250_U0_fifo_cout_drain_out_V_din_pass_1_q0 <= PE_wrapper250_U0_fifo_cout_drain_out_V_din_pass_1_out;
  end
  assign PE_wrapper250_U0_fifo_cout_drain_out_V_din_pass_1_in = PE_wrapper250_U0_fifo_cout_drain_out_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_PE_8_4_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_PE_8_4_V_full_n_pass_0_q0 <= fifo_cout_drain_PE_8_4_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_PE_8_4_V_full_n_pass_0_in = fifo_cout_drain_PE_8_4_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper250_U0_fifo_cout_drain_out_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper250_U0_fifo_cout_drain_out_V_write_pass_1_q0 <= PE_wrapper250_U0_fifo_cout_drain_out_V_write_pass_1_out;
  end
  assign PE_wrapper250_U0_fifo_cout_drain_out_V_write_pass_1_in = PE_wrapper250_U0_fifo_cout_drain_out_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper282_U0_fifo_cin_out_V_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper282_U0_fifo_cin_out_V_V_din_pass_1_q0 <= PE_wrapper282_U0_fifo_cin_out_V_V_din_pass_1_out;
  end
  assign PE_wrapper282_U0_fifo_cin_out_V_V_din_pass_1_in = PE_wrapper282_U0_fifo_cin_out_V_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_12_0_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_12_0_V_V_full_n_pass_0_q0 <= fifo_cin_PE_12_0_V_V_full_n_pass_0_out;
  end
  assign fifo_cin_PE_12_0_V_V_full_n_pass_0_in = fifo_cin_PE_12_0_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper282_U0_fifo_cin_out_V_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper282_U0_fifo_cin_out_V_V_write_pass_1_q0 <= PE_wrapper282_U0_fifo_cin_out_V_V_write_pass_1_out;
  end
  assign PE_wrapper282_U0_fifo_cin_out_V_V_write_pass_1_in = PE_wrapper282_U0_fifo_cin_out_V_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper237_U0_fifo_w_out_V_V_din_pass_2_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper237_U0_fifo_w_out_V_V_din_pass_2_q0 <= PE_wrapper237_U0_fifo_w_out_V_V_din_pass_2_out;
  end
  assign PE_wrapper237_U0_fifo_w_out_V_V_din_pass_2_in = PE_wrapper237_U0_fifo_w_out_V_V_din_pass_2_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_7_4_V_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_7_4_V_V_full_n_pass_1_q0 <= fifo_w_PE_7_4_V_V_full_n_pass_1_out;
  end
  assign fifo_w_PE_7_4_V_V_full_n_pass_1_in = fifo_w_PE_7_4_V_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper237_U0_fifo_w_out_V_V_write_pass_2_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper237_U0_fifo_w_out_V_V_write_pass_2_q0 <= PE_wrapper237_U0_fifo_w_out_V_V_write_pass_2_out;
  end
  assign PE_wrapper237_U0_fifo_w_out_V_V_write_pass_2_in = PE_wrapper237_U0_fifo_w_out_V_V_write_pass_2_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper283_U0_fifo_cin_out_V_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper283_U0_fifo_cin_out_V_V_din_pass_1_q0 <= PE_wrapper283_U0_fifo_cin_out_V_V_din_pass_1_out;
  end
  assign PE_wrapper283_U0_fifo_cin_out_V_V_din_pass_1_in = PE_wrapper283_U0_fifo_cin_out_V_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_12_1_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_12_1_V_V_full_n_pass_0_q0 <= fifo_cin_PE_12_1_V_V_full_n_pass_0_out;
  end
  assign fifo_cin_PE_12_1_V_V_full_n_pass_0_in = fifo_cin_PE_12_1_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper283_U0_fifo_cin_out_V_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper283_U0_fifo_cin_out_V_V_write_pass_1_q0 <= PE_wrapper283_U0_fifo_cin_out_V_V_write_pass_1_out;
  end
  assign PE_wrapper283_U0_fifo_cin_out_V_V_write_pass_1_in = PE_wrapper283_U0_fifo_cin_out_V_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper298_U0_fifo_w_out_V_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper298_U0_fifo_w_out_V_V_din_pass_1_q0 <= PE_wrapper298_U0_fifo_w_out_V_V_din_pass_1_out;
  end
  assign PE_wrapper298_U0_fifo_w_out_V_V_din_pass_1_in = PE_wrapper298_U0_fifo_w_out_V_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_12_5_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_12_5_V_V_full_n_pass_0_q0 <= fifo_w_PE_12_5_V_V_full_n_pass_0_out;
  end
  assign fifo_w_PE_12_5_V_V_full_n_pass_0_in = fifo_w_PE_12_5_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper298_U0_fifo_w_out_V_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper298_U0_fifo_w_out_V_V_write_pass_1_q0 <= PE_wrapper298_U0_fifo_w_out_V_V_write_pass_1_out;
  end
  assign PE_wrapper298_U0_fifo_w_out_V_V_write_pass_1_in = PE_wrapper298_U0_fifo_w_out_V_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper322_U0_fifo_w_out_V_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper322_U0_fifo_w_out_V_V_din_pass_1_q0 <= PE_wrapper322_U0_fifo_w_out_V_V_din_pass_1_out;
  end
  assign PE_wrapper322_U0_fifo_w_out_V_V_din_pass_1_in = PE_wrapper322_U0_fifo_w_out_V_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_14_5_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_14_5_V_V_full_n_pass_0_q0 <= fifo_w_PE_14_5_V_V_full_n_pass_0_out;
  end
  assign fifo_w_PE_14_5_V_V_full_n_pass_0_in = fifo_w_PE_14_5_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper322_U0_fifo_w_out_V_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper322_U0_fifo_w_out_V_V_write_pass_1_q0 <= PE_wrapper322_U0_fifo_w_out_V_V_write_pass_1_out;
  end
  assign PE_wrapper322_U0_fifo_w_out_V_V_write_pass_1_in = PE_wrapper322_U0_fifo_w_out_V_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper334_U0_fifo_w_out_V_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper334_U0_fifo_w_out_V_V_din_pass_1_q0 <= PE_wrapper334_U0_fifo_w_out_V_V_din_pass_1_out;
  end
  assign PE_wrapper334_U0_fifo_w_out_V_V_din_pass_1_in = PE_wrapper334_U0_fifo_w_out_V_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_15_5_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_15_5_V_V_full_n_pass_0_q0 <= fifo_w_PE_15_5_V_V_full_n_pass_0_out;
  end
  assign fifo_w_PE_15_5_V_V_full_n_pass_0_in = fifo_w_PE_15_5_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper334_U0_fifo_w_out_V_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper334_U0_fifo_w_out_V_V_write_pass_1_q0 <= PE_wrapper334_U0_fifo_w_out_V_V_write_pass_1_out;
  end
  assign PE_wrapper334_U0_fifo_w_out_V_V_write_pass_1_in = PE_wrapper334_U0_fifo_w_out_V_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_cout_drain_IO_L1_out_1_13_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_cout_drain_IO_L1_out_1_13_V_V_full_n_pass_0_q0 <= fifo_cout_drain_cout_drain_IO_L1_out_1_13_V_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_cout_drain_IO_L1_out_1_13_V_V_full_n_pass_0_in = fifo_cout_drain_cout_drain_IO_L1_out_1_13_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper309_U0_fifo_cin_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper309_U0_fifo_cin_out_V_V_din_pass_0_q0 <= PE_wrapper309_U0_fifo_cin_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper309_U0_fifo_cin_out_V_V_din_pass_0_in = PE_wrapper309_U0_fifo_cin_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper309_U0_fifo_cin_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper309_U0_fifo_cin_out_V_V_write_pass_0_q0 <= PE_wrapper309_U0_fifo_cin_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper309_U0_fifo_cin_out_V_V_write_pass_0_in = PE_wrapper309_U0_fifo_cin_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_9_4_V_V_full_n_pass_2_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_9_4_V_V_full_n_pass_2_q0 <= fifo_w_PE_9_4_V_V_full_n_pass_2_out;
  end
  assign fifo_w_PE_9_4_V_V_full_n_pass_2_in = fifo_w_PE_9_4_V_V_full_n_pass_2_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper333_U0_fifo_w_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper333_U0_fifo_w_out_V_V_din_pass_0_q0 <= PE_wrapper333_U0_fifo_w_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper333_U0_fifo_w_out_V_V_din_pass_0_in = PE_wrapper333_U0_fifo_w_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper333_U0_fifo_w_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper333_U0_fifo_w_out_V_V_write_pass_0_q0 <= PE_wrapper333_U0_fifo_w_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper333_U0_fifo_w_out_V_V_write_pass_0_in = PE_wrapper333_U0_fifo_w_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [63:0] cout_drain_IO_L1_out_wrapper440_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper440_U0_fifo_cout_drain_out_V_V_din_pass_0_q0 <= cout_drain_IO_L1_out_wrapper440_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper440_U0_fifo_cout_drain_out_V_V_din_pass_0_in = cout_drain_IO_L1_out_wrapper440_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  cout_drain_IO_L1_out_wrapper440_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper440_U0_fifo_cout_drain_out_V_V_write_pass_0_q0 <= cout_drain_IO_L1_out_wrapper440_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper440_U0_fifo_cout_drain_out_V_V_write_pass_0_in = cout_drain_IO_L1_out_wrapper440_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_9_4_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_9_4_V_V_full_n_pass_0_q0 <= fifo_cin_PE_9_4_V_V_full_n_pass_0_out;
  end
  assign fifo_cin_PE_9_4_V_V_full_n_pass_0_in = fifo_cin_PE_9_4_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_PE_11_4_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_PE_11_4_V_full_n_pass_1_q0 <= fifo_cout_drain_PE_11_4_V_full_n_pass_1_out;
  end
  assign fifo_cout_drain_PE_11_4_V_full_n_pass_1_in = fifo_cout_drain_PE_11_4_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_cout_drain_IO_L1_out_4_7_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_cout_drain_IO_L1_out_4_7_V_V_full_n_pass_0_q0 <= fifo_cout_drain_cout_drain_IO_L1_out_4_7_V_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_cout_drain_IO_L1_out_4_7_V_V_full_n_pass_0_in = fifo_cout_drain_cout_drain_IO_L1_out_4_7_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg [31:0] PE_wrapper306_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper306_U0_fifo_cout_drain_out_V_din_pass_0_q0 <= PE_wrapper306_U0_fifo_cout_drain_out_V_din_pass_0_out;
  end
  assign PE_wrapper306_U0_fifo_cout_drain_out_V_din_pass_0_in = PE_wrapper306_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper306_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper306_U0_fifo_cout_drain_out_V_write_pass_0_q0 <= PE_wrapper306_U0_fifo_cout_drain_out_V_write_pass_0_out;
  end
  assign PE_wrapper306_U0_fifo_cout_drain_out_V_write_pass_0_in = PE_wrapper306_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_12_2_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_12_2_V_V_full_n_pass_0_q0 <= fifo_w_PE_12_2_V_V_full_n_pass_0_out;
  end
  assign fifo_w_PE_12_2_V_V_full_n_pass_0_in = fifo_w_PE_12_2_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_PE_6_4_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_PE_6_4_V_full_n_pass_1_q0 <= fifo_cout_drain_PE_6_4_V_full_n_pass_1_out;
  end
  assign fifo_cout_drain_PE_6_4_V_full_n_pass_1_in = fifo_cout_drain_PE_6_4_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_15_2_V_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_15_2_V_V_full_n_pass_1_q0 <= fifo_cin_PE_15_2_V_V_full_n_pass_1_out;
  end
  assign fifo_cin_PE_15_2_V_V_full_n_pass_1_in = fifo_cin_PE_15_2_V_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper309_U0_fifo_w_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper309_U0_fifo_w_out_V_V_din_pass_0_q0 <= PE_wrapper309_U0_fifo_w_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper309_U0_fifo_w_out_V_V_din_pass_0_in = PE_wrapper309_U0_fifo_w_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper309_U0_fifo_w_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper309_U0_fifo_w_out_V_V_write_pass_0_q0 <= PE_wrapper309_U0_fifo_w_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper309_U0_fifo_w_out_V_V_write_pass_0_in = PE_wrapper309_U0_fifo_w_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_15_2_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_15_2_V_V_full_n_pass_0_q0 <= fifo_w_PE_15_2_V_V_full_n_pass_0_out;
  end
  assign fifo_w_PE_15_2_V_V_full_n_pass_0_in = fifo_w_PE_15_2_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg [63:0] cout_drain_IO_L1_out_wrapper418_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper418_U0_fifo_cout_drain_out_V_V_din_pass_0_q0 <= cout_drain_IO_L1_out_wrapper418_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper418_U0_fifo_cout_drain_out_V_V_din_pass_0_in = cout_drain_IO_L1_out_wrapper418_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  cout_drain_IO_L1_out_wrapper418_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper418_U0_fifo_cout_drain_out_V_V_write_pass_0_q0 <= cout_drain_IO_L1_out_wrapper418_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper418_U0_fifo_cout_drain_out_V_V_write_pass_0_in = cout_drain_IO_L1_out_wrapper418_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_cout_drain_IO_L1_out_3_13_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_cout_drain_IO_L1_out_3_13_V_V_full_n_pass_0_q0 <= fifo_cout_drain_cout_drain_IO_L1_out_3_13_V_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_cout_drain_IO_L1_out_3_13_V_V_full_n_pass_0_in = fifo_cout_drain_cout_drain_IO_L1_out_3_13_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] w_IO_L2_in147_U0_fifo_w_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    w_IO_L2_in147_U0_fifo_w_out_V_V_din_pass_0_q0 <= w_IO_L2_in147_U0_fifo_w_out_V_V_din_pass_0_out;
  end
  assign w_IO_L2_in147_U0_fifo_w_out_V_V_din_pass_0_in = w_IO_L2_in147_U0_fifo_w_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  w_IO_L2_in147_U0_fifo_w_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    w_IO_L2_in147_U0_fifo_w_out_V_V_write_pass_0_q0 <= w_IO_L2_in147_U0_fifo_w_out_V_V_write_pass_0_out;
  end
  assign w_IO_L2_in147_U0_fifo_w_out_V_V_write_pass_0_in = w_IO_L2_in147_U0_fifo_w_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_w_w_IO_L2_in_12_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_w_IO_L2_in_12_V_V_full_n_pass_0_q0 <= fifo_w_w_IO_L2_in_12_V_V_full_n_pass_0_out;
  end
  assign fifo_w_w_IO_L2_in_12_V_V_full_n_pass_0_in = fifo_w_w_IO_L2_in_12_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_13_3_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_13_3_V_V_full_n_pass_0_q0 <= fifo_cin_PE_13_3_V_V_full_n_pass_0_out;
  end
  assign fifo_cin_PE_13_3_V_V_full_n_pass_0_in = fifo_cin_PE_13_3_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper285_U0_fifo_w_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper285_U0_fifo_w_out_V_V_din_pass_0_q0 <= PE_wrapper285_U0_fifo_w_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper285_U0_fifo_w_out_V_V_din_pass_0_in = PE_wrapper285_U0_fifo_w_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper285_U0_fifo_w_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper285_U0_fifo_w_out_V_V_write_pass_0_q0 <= PE_wrapper285_U0_fifo_w_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper285_U0_fifo_w_out_V_V_write_pass_0_in = PE_wrapper285_U0_fifo_w_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper306_U0_fifo_w_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper306_U0_fifo_w_out_V_V_din_pass_0_q0 <= PE_wrapper306_U0_fifo_w_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper306_U0_fifo_w_out_V_V_din_pass_0_in = PE_wrapper306_U0_fifo_w_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper306_U0_fifo_w_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper306_U0_fifo_w_out_V_V_write_pass_0_q0 <= PE_wrapper306_U0_fifo_w_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper306_U0_fifo_w_out_V_V_write_pass_0_in = PE_wrapper306_U0_fifo_w_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [31:0] PE_wrapper333_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper333_U0_fifo_cout_drain_out_V_din_pass_0_q0 <= PE_wrapper333_U0_fifo_cout_drain_out_V_din_pass_0_out;
  end
  assign PE_wrapper333_U0_fifo_cout_drain_out_V_din_pass_0_in = PE_wrapper333_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper333_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper333_U0_fifo_cout_drain_out_V_write_pass_0_q0 <= PE_wrapper333_U0_fifo_cout_drain_out_V_write_pass_0_out;
  end
  assign PE_wrapper333_U0_fifo_cout_drain_out_V_write_pass_0_in = PE_wrapper333_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [63:0] cout_drain_IO_L1_out_wrapper386_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper386_U0_fifo_cout_drain_out_V_V_din_pass_0_q0 <= cout_drain_IO_L1_out_wrapper386_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper386_U0_fifo_cout_drain_out_V_V_din_pass_0_in = cout_drain_IO_L1_out_wrapper386_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  cout_drain_IO_L1_out_wrapper386_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper386_U0_fifo_cout_drain_out_V_V_write_pass_0_q0 <= cout_drain_IO_L1_out_wrapper386_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper386_U0_fifo_cout_drain_out_V_V_write_pass_0_in = cout_drain_IO_L1_out_wrapper386_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper262_U0_fifo_w_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper262_U0_fifo_w_out_V_V_din_pass_0_q0 <= PE_wrapper262_U0_fifo_w_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper262_U0_fifo_w_out_V_V_din_pass_0_in = PE_wrapper262_U0_fifo_w_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper262_U0_fifo_w_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper262_U0_fifo_w_out_V_V_write_pass_0_q0 <= PE_wrapper262_U0_fifo_w_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper262_U0_fifo_w_out_V_V_write_pass_0_in = PE_wrapper262_U0_fifo_w_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper306_U0_fifo_cin_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper306_U0_fifo_cin_out_V_V_din_pass_0_q0 <= PE_wrapper306_U0_fifo_cin_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper306_U0_fifo_cin_out_V_V_din_pass_0_in = PE_wrapper306_U0_fifo_cin_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper306_U0_fifo_cin_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper306_U0_fifo_cin_out_V_V_write_pass_0_q0 <= PE_wrapper306_U0_fifo_cin_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper306_U0_fifo_cin_out_V_V_write_pass_0_in = PE_wrapper306_U0_fifo_cin_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_11_3_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_11_3_V_V_full_n_pass_0_q0 <= fifo_cin_PE_11_3_V_V_full_n_pass_0_out;
  end
  assign fifo_cin_PE_11_3_V_V_full_n_pass_0_in = fifo_cin_PE_11_3_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_15_3_V_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_15_3_V_V_full_n_pass_1_q0 <= fifo_cin_PE_15_3_V_V_full_n_pass_1_out;
  end
  assign fifo_cin_PE_15_3_V_V_full_n_pass_1_in = fifo_cin_PE_15_3_V_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_PE_12_1_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_PE_12_1_V_full_n_pass_0_q0 <= fifo_cout_drain_PE_12_1_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_PE_12_1_V_full_n_pass_0_in = fifo_cout_drain_PE_12_1_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg [31:0] PE_wrapper285_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper285_U0_fifo_cout_drain_out_V_din_pass_0_q0 <= PE_wrapper285_U0_fifo_cout_drain_out_V_din_pass_0_out;
  end
  assign PE_wrapper285_U0_fifo_cout_drain_out_V_din_pass_0_in = PE_wrapper285_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper285_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper285_U0_fifo_cout_drain_out_V_write_pass_0_q0 <= PE_wrapper285_U0_fifo_cout_drain_out_V_write_pass_0_out;
  end
  assign PE_wrapper285_U0_fifo_cout_drain_out_V_write_pass_0_in = PE_wrapper285_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_13_0_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_13_0_V_V_full_n_pass_0_q0 <= fifo_cin_PE_13_0_V_V_full_n_pass_0_out;
  end
  assign fifo_cin_PE_13_0_V_V_full_n_pass_0_in = fifo_cin_PE_13_0_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] w_IO_L2_in147_U0_fifo_w_local_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    w_IO_L2_in147_U0_fifo_w_local_out_V_V_din_pass_0_q0 <= w_IO_L2_in147_U0_fifo_w_local_out_V_V_din_pass_0_out;
  end
  assign w_IO_L2_in147_U0_fifo_w_local_out_V_V_din_pass_0_in = w_IO_L2_in147_U0_fifo_w_local_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  w_IO_L2_in147_U0_fifo_w_local_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    w_IO_L2_in147_U0_fifo_w_local_out_V_V_write_pass_0_q0 <= w_IO_L2_in147_U0_fifo_w_local_out_V_V_write_pass_0_out;
  end
  assign w_IO_L2_in147_U0_fifo_w_local_out_V_V_write_pass_0_in = w_IO_L2_in147_U0_fifo_w_local_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [63:0] cout_drain_IO_L1_out_wrapper437_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper437_U0_fifo_cout_drain_out_V_V_din_pass_0_q0 <= cout_drain_IO_L1_out_wrapper437_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper437_U0_fifo_cout_drain_out_V_V_din_pass_0_in = cout_drain_IO_L1_out_wrapper437_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  cout_drain_IO_L1_out_wrapper437_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper437_U0_fifo_cout_drain_out_V_V_write_pass_0_q0 <= cout_drain_IO_L1_out_wrapper437_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper437_U0_fifo_cout_drain_out_V_V_write_pass_0_in = cout_drain_IO_L1_out_wrapper437_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_PE_12_3_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_PE_12_3_V_full_n_pass_0_q0 <= fifo_cout_drain_PE_12_3_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_PE_12_3_V_full_n_pass_0_in = fifo_cout_drain_PE_12_3_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_13_3_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_13_3_V_V_full_n_pass_0_q0 <= fifo_w_PE_13_3_V_V_full_n_pass_0_out;
  end
  assign fifo_w_PE_13_3_V_V_full_n_pass_0_in = fifo_w_PE_13_3_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper296_U0_fifo_cin_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper296_U0_fifo_cin_out_V_V_din_pass_0_q0 <= PE_wrapper296_U0_fifo_cin_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper296_U0_fifo_cin_out_V_V_din_pass_0_in = PE_wrapper296_U0_fifo_cin_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper296_U0_fifo_cin_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper296_U0_fifo_cin_out_V_V_write_pass_0_q0 <= PE_wrapper296_U0_fifo_cin_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper296_U0_fifo_cin_out_V_V_write_pass_0_in = PE_wrapper296_U0_fifo_cin_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_11_3_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_11_3_V_V_full_n_pass_0_q0 <= fifo_w_PE_11_3_V_V_full_n_pass_0_out;
  end
  assign fifo_w_PE_11_3_V_V_full_n_pass_0_in = fifo_w_PE_11_3_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper296_U0_fifo_w_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper296_U0_fifo_w_out_V_V_din_pass_0_q0 <= PE_wrapper296_U0_fifo_w_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper296_U0_fifo_w_out_V_V_din_pass_0_in = PE_wrapper296_U0_fifo_w_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper296_U0_fifo_w_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper296_U0_fifo_w_out_V_V_write_pass_0_q0 <= PE_wrapper296_U0_fifo_w_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper296_U0_fifo_w_out_V_V_write_pass_0_in = PE_wrapper296_U0_fifo_w_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [31:0] PE_wrapper296_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper296_U0_fifo_cout_drain_out_V_din_pass_0_q0 <= PE_wrapper296_U0_fifo_cout_drain_out_V_din_pass_0_out;
  end
  assign PE_wrapper296_U0_fifo_cout_drain_out_V_din_pass_0_in = PE_wrapper296_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper296_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper296_U0_fifo_cout_drain_out_V_write_pass_0_q0 <= PE_wrapper296_U0_fifo_cout_drain_out_V_write_pass_0_out;
  end
  assign PE_wrapper296_U0_fifo_cout_drain_out_V_write_pass_0_in = PE_wrapper296_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper262_U0_fifo_cin_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper262_U0_fifo_cin_out_V_V_din_pass_0_q0 <= PE_wrapper262_U0_fifo_cin_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper262_U0_fifo_cin_out_V_V_din_pass_0_in = PE_wrapper262_U0_fifo_cin_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper262_U0_fifo_cin_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper262_U0_fifo_cin_out_V_V_write_pass_0_q0 <= PE_wrapper262_U0_fifo_cin_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper262_U0_fifo_cin_out_V_V_write_pass_0_in = PE_wrapper262_U0_fifo_cin_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_PE_10_4_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_PE_10_4_V_full_n_pass_1_q0 <= fifo_cout_drain_PE_10_4_V_full_n_pass_1_out;
  end
  assign fifo_cout_drain_PE_10_4_V_full_n_pass_1_in = fifo_cout_drain_PE_10_4_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_13_0_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_13_0_V_V_full_n_pass_0_q0 <= fifo_w_PE_13_0_V_V_full_n_pass_0_out;
  end
  assign fifo_w_PE_13_0_V_V_full_n_pass_0_in = fifo_w_PE_13_0_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg [63:0] cout_drain_IO_L1_out_boundary_wrapper399_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_boundary_wrapper399_U0_fifo_cout_drain_out_V_V_din_pass_0_q0 <= cout_drain_IO_L1_out_boundary_wrapper399_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  end
  assign cout_drain_IO_L1_out_boundary_wrapper399_U0_fifo_cout_drain_out_V_V_din_pass_0_in = cout_drain_IO_L1_out_boundary_wrapper399_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  cout_drain_IO_L1_out_boundary_wrapper399_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_boundary_wrapper399_U0_fifo_cout_drain_out_V_V_write_pass_0_q0 <= cout_drain_IO_L1_out_boundary_wrapper399_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  end
  assign cout_drain_IO_L1_out_boundary_wrapper399_U0_fifo_cout_drain_out_V_V_write_pass_0_in = cout_drain_IO_L1_out_boundary_wrapper399_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_12_2_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_12_2_V_V_full_n_pass_0_q0 <= fifo_cin_PE_12_2_V_V_full_n_pass_0_out;
  end
  assign fifo_cin_PE_12_2_V_V_full_n_pass_0_in = fifo_cin_PE_12_2_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_cout_drain_IO_L1_out_4_12_V_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_cout_drain_IO_L1_out_4_12_V_V_full_n_pass_1_q0 <= fifo_cout_drain_cout_drain_IO_L1_out_4_12_V_V_full_n_pass_1_out;
  end
  assign fifo_cout_drain_cout_drain_IO_L1_out_4_12_V_V_full_n_pass_1_in = fifo_cout_drain_cout_drain_IO_L1_out_4_12_V_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper285_U0_fifo_cin_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper285_U0_fifo_cin_out_V_V_din_pass_0_q0 <= PE_wrapper285_U0_fifo_cin_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper285_U0_fifo_cin_out_V_V_din_pass_0_in = PE_wrapper285_U0_fifo_cin_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper285_U0_fifo_cin_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper285_U0_fifo_cin_out_V_V_write_pass_0_q0 <= PE_wrapper285_U0_fifo_cin_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper285_U0_fifo_cin_out_V_V_write_pass_0_in = PE_wrapper285_U0_fifo_cin_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [31:0] PE_wrapper309_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper309_U0_fifo_cout_drain_out_V_din_pass_0_q0 <= PE_wrapper309_U0_fifo_cout_drain_out_V_din_pass_0_out;
  end
  assign PE_wrapper309_U0_fifo_cout_drain_out_V_din_pass_0_in = PE_wrapper309_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper309_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper309_U0_fifo_cout_drain_out_V_write_pass_0_q0 <= PE_wrapper309_U0_fifo_cout_drain_out_V_write_pass_0_out;
  end
  assign PE_wrapper309_U0_fifo_cout_drain_out_V_write_pass_0_in = PE_wrapper309_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  ap_done_Boundary_X0Y4_To_X2Y4_q0;
  always @ (posedge ap_clk) begin
    ap_done_Boundary_X0Y4_To_X2Y4_q0 <= ap_done_Boundary_X0Y4_To_X2Y4_out;
  end
  assign ap_done_Boundary_X0Y4_To_X2Y4_in = ap_done_Boundary_X0Y4_To_X2Y4_q0;
  (* dont_touch = "yes" *) reg  ap_start_Boundary_X0Y6_To_X2Y6_q0;
  always @ (posedge ap_clk) begin
    ap_start_Boundary_X0Y6_To_X2Y6_q0 <= ap_start_Boundary_X0Y6_To_X2Y6_out;
  end
  assign ap_start_Boundary_X0Y6_To_X2Y6_in = ap_start_Boundary_X0Y6_To_X2Y6_q0;
  (* dont_touch = "yes" *) reg  ap_rst_n_Boundary_X0Y6_To_X2Y6_q0;
  always @ (posedge ap_clk) begin
    ap_rst_n_Boundary_X0Y6_To_X2Y6_q0 <= ap_rst_n_Boundary_X0Y6_To_X2Y6_out;
  end
  assign ap_rst_n_Boundary_X0Y6_To_X2Y6_in = ap_rst_n_Boundary_X0Y6_To_X2Y6_q0;
  (* dont_touch = "yes" *) reg [63:0] cout_drain_IO_L1_out_wrapper402_U0_fifo_cout_drain_out_V_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper402_U0_fifo_cout_drain_out_V_V_din_pass_1_q0 <= cout_drain_IO_L1_out_wrapper402_U0_fifo_cout_drain_out_V_V_din_pass_1_out;
  end
  assign cout_drain_IO_L1_out_wrapper402_U0_fifo_cout_drain_out_V_V_din_pass_1_in = cout_drain_IO_L1_out_wrapper402_U0_fifo_cout_drain_out_V_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_cout_drain_IO_L1_out_2_12_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_cout_drain_IO_L1_out_2_12_V_V_full_n_pass_0_q0 <= fifo_cout_drain_cout_drain_IO_L1_out_2_12_V_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_cout_drain_IO_L1_out_2_12_V_V_full_n_pass_0_in = fifo_cout_drain_cout_drain_IO_L1_out_2_12_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  cout_drain_IO_L1_out_wrapper402_U0_fifo_cout_drain_out_V_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper402_U0_fifo_cout_drain_out_V_V_write_pass_1_q0 <= cout_drain_IO_L1_out_wrapper402_U0_fifo_cout_drain_out_V_V_write_pass_1_out;
  end
  assign cout_drain_IO_L1_out_wrapper402_U0_fifo_cout_drain_out_V_V_write_pass_1_in = cout_drain_IO_L1_out_wrapper402_U0_fifo_cout_drain_out_V_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [31:0] PE_wrapper286_U0_fifo_cout_drain_out_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper286_U0_fifo_cout_drain_out_V_din_pass_1_q0 <= PE_wrapper286_U0_fifo_cout_drain_out_V_din_pass_1_out;
  end
  assign PE_wrapper286_U0_fifo_cout_drain_out_V_din_pass_1_in = PE_wrapper286_U0_fifo_cout_drain_out_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_PE_11_4_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_PE_11_4_V_full_n_pass_0_q0 <= fifo_cout_drain_PE_11_4_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_PE_11_4_V_full_n_pass_0_in = fifo_cout_drain_PE_11_4_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper286_U0_fifo_cout_drain_out_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper286_U0_fifo_cout_drain_out_V_write_pass_1_q0 <= PE_wrapper286_U0_fifo_cout_drain_out_V_write_pass_1_out;
  end
  assign PE_wrapper286_U0_fifo_cout_drain_out_V_write_pass_1_in = PE_wrapper286_U0_fifo_cout_drain_out_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [31:0] PE_wrapper226_U0_fifo_cout_drain_out_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper226_U0_fifo_cout_drain_out_V_din_pass_1_q0 <= PE_wrapper226_U0_fifo_cout_drain_out_V_din_pass_1_out;
  end
  assign PE_wrapper226_U0_fifo_cout_drain_out_V_din_pass_1_in = PE_wrapper226_U0_fifo_cout_drain_out_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_PE_6_4_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_PE_6_4_V_full_n_pass_0_q0 <= fifo_cout_drain_PE_6_4_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_PE_6_4_V_full_n_pass_0_in = fifo_cout_drain_PE_6_4_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper226_U0_fifo_cout_drain_out_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper226_U0_fifo_cout_drain_out_V_write_pass_1_q0 <= PE_wrapper226_U0_fifo_cout_drain_out_V_write_pass_1_out;
  end
  assign PE_wrapper226_U0_fifo_cout_drain_out_V_write_pass_1_in = PE_wrapper226_U0_fifo_cout_drain_out_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper320_U0_fifo_cin_out_V_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper320_U0_fifo_cin_out_V_V_din_pass_1_q0 <= PE_wrapper320_U0_fifo_cin_out_V_V_din_pass_1_out;
  end
  assign PE_wrapper320_U0_fifo_cin_out_V_V_din_pass_1_in = PE_wrapper320_U0_fifo_cin_out_V_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_15_2_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_15_2_V_V_full_n_pass_0_q0 <= fifo_cin_PE_15_2_V_V_full_n_pass_0_out;
  end
  assign fifo_cin_PE_15_2_V_V_full_n_pass_0_in = fifo_cin_PE_15_2_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper320_U0_fifo_cin_out_V_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper320_U0_fifo_cin_out_V_V_write_pass_1_q0 <= PE_wrapper320_U0_fifo_cin_out_V_V_write_pass_1_out;
  end
  assign PE_wrapper320_U0_fifo_cin_out_V_V_write_pass_1_in = PE_wrapper320_U0_fifo_cin_out_V_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper321_U0_fifo_cin_out_V_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper321_U0_fifo_cin_out_V_V_din_pass_1_q0 <= PE_wrapper321_U0_fifo_cin_out_V_V_din_pass_1_out;
  end
  assign PE_wrapper321_U0_fifo_cin_out_V_V_din_pass_1_in = PE_wrapper321_U0_fifo_cin_out_V_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_15_3_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_15_3_V_V_full_n_pass_0_q0 <= fifo_cin_PE_15_3_V_V_full_n_pass_0_out;
  end
  assign fifo_cin_PE_15_3_V_V_full_n_pass_0_in = fifo_cin_PE_15_3_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper321_U0_fifo_cin_out_V_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper321_U0_fifo_cin_out_V_V_write_pass_1_q0 <= PE_wrapper321_U0_fifo_cin_out_V_V_write_pass_1_out;
  end
  assign PE_wrapper321_U0_fifo_cin_out_V_V_write_pass_1_in = PE_wrapper321_U0_fifo_cin_out_V_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [31:0] PE_wrapper274_U0_fifo_cout_drain_out_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper274_U0_fifo_cout_drain_out_V_din_pass_1_q0 <= PE_wrapper274_U0_fifo_cout_drain_out_V_din_pass_1_out;
  end
  assign PE_wrapper274_U0_fifo_cout_drain_out_V_din_pass_1_in = PE_wrapper274_U0_fifo_cout_drain_out_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_PE_10_4_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_PE_10_4_V_full_n_pass_0_q0 <= fifo_cout_drain_PE_10_4_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_PE_10_4_V_full_n_pass_0_in = fifo_cout_drain_PE_10_4_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper274_U0_fifo_cout_drain_out_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper274_U0_fifo_cout_drain_out_V_write_pass_1_q0 <= PE_wrapper274_U0_fifo_cout_drain_out_V_write_pass_1_out;
  end
  assign PE_wrapper274_U0_fifo_cout_drain_out_V_write_pass_1_in = PE_wrapper274_U0_fifo_cout_drain_out_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [63:0] cout_drain_IO_L1_out_wrapper434_U0_fifo_cout_drain_out_V_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper434_U0_fifo_cout_drain_out_V_V_din_pass_1_q0 <= cout_drain_IO_L1_out_wrapper434_U0_fifo_cout_drain_out_V_V_din_pass_1_out;
  end
  assign cout_drain_IO_L1_out_wrapper434_U0_fifo_cout_drain_out_V_V_din_pass_1_in = cout_drain_IO_L1_out_wrapper434_U0_fifo_cout_drain_out_V_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_cout_drain_IO_L1_out_4_12_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_cout_drain_IO_L1_out_4_12_V_V_full_n_pass_0_q0 <= fifo_cout_drain_cout_drain_IO_L1_out_4_12_V_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_cout_drain_IO_L1_out_4_12_V_V_full_n_pass_0_in = fifo_cout_drain_cout_drain_IO_L1_out_4_12_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  cout_drain_IO_L1_out_wrapper434_U0_fifo_cout_drain_out_V_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper434_U0_fifo_cout_drain_out_V_V_write_pass_1_q0 <= cout_drain_IO_L1_out_wrapper434_U0_fifo_cout_drain_out_V_V_write_pass_1_out;
  end
  assign cout_drain_IO_L1_out_wrapper434_U0_fifo_cout_drain_out_V_V_write_pass_1_in = cout_drain_IO_L1_out_wrapper434_U0_fifo_cout_drain_out_V_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper262_U0_fifo_w_out_V_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper262_U0_fifo_w_out_V_V_din_pass_1_q0 <= PE_wrapper262_U0_fifo_w_out_V_V_din_pass_1_out;
  end
  assign PE_wrapper262_U0_fifo_w_out_V_V_din_pass_1_in = PE_wrapper262_U0_fifo_w_out_V_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_9_5_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_9_5_V_V_full_n_pass_0_q0 <= fifo_w_PE_9_5_V_V_full_n_pass_0_out;
  end
  assign fifo_w_PE_9_5_V_V_full_n_pass_0_in = fifo_w_PE_9_5_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper262_U0_fifo_w_out_V_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper262_U0_fifo_w_out_V_V_write_pass_1_q0 <= PE_wrapper262_U0_fifo_w_out_V_V_write_pass_1_out;
  end
  assign PE_wrapper262_U0_fifo_w_out_V_V_write_pass_1_in = PE_wrapper262_U0_fifo_w_out_V_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper298_U0_fifo_w_out_V_V_din_pass_2_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper298_U0_fifo_w_out_V_V_din_pass_2_q0 <= PE_wrapper298_U0_fifo_w_out_V_V_din_pass_2_out;
  end
  assign PE_wrapper298_U0_fifo_w_out_V_V_din_pass_2_in = PE_wrapper298_U0_fifo_w_out_V_V_din_pass_2_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_12_5_V_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_12_5_V_V_full_n_pass_1_q0 <= fifo_w_PE_12_5_V_V_full_n_pass_1_out;
  end
  assign fifo_w_PE_12_5_V_V_full_n_pass_1_in = fifo_w_PE_12_5_V_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper298_U0_fifo_w_out_V_V_write_pass_2_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper298_U0_fifo_w_out_V_V_write_pass_2_q0 <= PE_wrapper298_U0_fifo_w_out_V_V_write_pass_2_out;
  end
  assign PE_wrapper298_U0_fifo_w_out_V_V_write_pass_2_in = PE_wrapper298_U0_fifo_w_out_V_V_write_pass_2_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper322_U0_fifo_w_out_V_V_din_pass_2_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper322_U0_fifo_w_out_V_V_din_pass_2_q0 <= PE_wrapper322_U0_fifo_w_out_V_V_din_pass_2_out;
  end
  assign PE_wrapper322_U0_fifo_w_out_V_V_din_pass_2_in = PE_wrapper322_U0_fifo_w_out_V_V_din_pass_2_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_14_5_V_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_14_5_V_V_full_n_pass_1_q0 <= fifo_w_PE_14_5_V_V_full_n_pass_1_out;
  end
  assign fifo_w_PE_14_5_V_V_full_n_pass_1_in = fifo_w_PE_14_5_V_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper322_U0_fifo_w_out_V_V_write_pass_2_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper322_U0_fifo_w_out_V_V_write_pass_2_q0 <= PE_wrapper322_U0_fifo_w_out_V_V_write_pass_2_out;
  end
  assign PE_wrapper322_U0_fifo_w_out_V_V_write_pass_2_in = PE_wrapper322_U0_fifo_w_out_V_V_write_pass_2_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper334_U0_fifo_w_out_V_V_din_pass_2_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper334_U0_fifo_w_out_V_V_din_pass_2_q0 <= PE_wrapper334_U0_fifo_w_out_V_V_din_pass_2_out;
  end
  assign PE_wrapper334_U0_fifo_w_out_V_V_din_pass_2_in = PE_wrapper334_U0_fifo_w_out_V_V_din_pass_2_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_15_5_V_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_15_5_V_V_full_n_pass_1_q0 <= fifo_w_PE_15_5_V_V_full_n_pass_1_out;
  end
  assign fifo_w_PE_15_5_V_V_full_n_pass_1_in = fifo_w_PE_15_5_V_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper334_U0_fifo_w_out_V_V_write_pass_2_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper334_U0_fifo_w_out_V_V_write_pass_2_q0 <= PE_wrapper334_U0_fifo_w_out_V_V_write_pass_2_out;
  end
  assign PE_wrapper334_U0_fifo_w_out_V_V_write_pass_2_in = PE_wrapper334_U0_fifo_w_out_V_V_write_pass_2_q0;
  (* dont_touch = "yes" *) reg [63:0] cout_drain_IO_L1_out_wrapper385_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper385_U0_fifo_cout_drain_out_V_V_din_pass_0_q0 <= cout_drain_IO_L1_out_wrapper385_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper385_U0_fifo_cout_drain_out_V_V_din_pass_0_in = cout_drain_IO_L1_out_wrapper385_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  cout_drain_IO_L1_out_wrapper385_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper385_U0_fifo_cout_drain_out_V_V_write_pass_0_q0 <= cout_drain_IO_L1_out_wrapper385_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper385_U0_fifo_cout_drain_out_V_V_write_pass_0_in = cout_drain_IO_L1_out_wrapper385_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_13_4_V_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_13_4_V_V_full_n_pass_1_q0 <= fifo_cin_PE_13_4_V_V_full_n_pass_1_out;
  end
  assign fifo_cin_PE_13_4_V_V_full_n_pass_1_in = fifo_cin_PE_13_4_V_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_PE_8_4_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_PE_8_4_V_full_n_pass_1_q0 <= fifo_cout_drain_PE_8_4_V_full_n_pass_1_out;
  end
  assign fifo_cout_drain_PE_8_4_V_full_n_pass_1_in = fifo_cout_drain_PE_8_4_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper310_U0_fifo_w_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper310_U0_fifo_w_out_V_V_din_pass_0_q0 <= PE_wrapper310_U0_fifo_w_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper310_U0_fifo_w_out_V_V_din_pass_0_in = PE_wrapper310_U0_fifo_w_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper310_U0_fifo_w_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper310_U0_fifo_w_out_V_V_write_pass_0_q0 <= PE_wrapper310_U0_fifo_w_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper310_U0_fifo_w_out_V_V_write_pass_0_in = PE_wrapper310_U0_fifo_w_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [63:0] cout_drain_IO_L1_out_wrapper439_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper439_U0_fifo_cout_drain_out_V_V_din_pass_0_q0 <= cout_drain_IO_L1_out_wrapper439_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper439_U0_fifo_cout_drain_out_V_V_din_pass_0_in = cout_drain_IO_L1_out_wrapper439_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  cout_drain_IO_L1_out_wrapper439_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper439_U0_fifo_cout_drain_out_V_V_write_pass_0_q0 <= cout_drain_IO_L1_out_wrapper439_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper439_U0_fifo_cout_drain_out_V_V_write_pass_0_in = cout_drain_IO_L1_out_wrapper439_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [31:0] PE_wrapper310_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper310_U0_fifo_cout_drain_out_V_din_pass_0_q0 <= PE_wrapper310_U0_fifo_cout_drain_out_V_din_pass_0_out;
  end
  assign PE_wrapper310_U0_fifo_cout_drain_out_V_din_pass_0_in = PE_wrapper310_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper310_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper310_U0_fifo_cout_drain_out_V_write_pass_0_q0 <= PE_wrapper310_U0_fifo_cout_drain_out_V_write_pass_0_out;
  end
  assign PE_wrapper310_U0_fifo_cout_drain_out_V_write_pass_0_in = PE_wrapper310_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper295_U0_fifo_w_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper295_U0_fifo_w_out_V_V_din_pass_0_q0 <= PE_wrapper295_U0_fifo_w_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper295_U0_fifo_w_out_V_V_din_pass_0_in = PE_wrapper295_U0_fifo_w_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper295_U0_fifo_w_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper295_U0_fifo_w_out_V_V_write_pass_0_q0 <= PE_wrapper295_U0_fifo_w_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper295_U0_fifo_w_out_V_V_write_pass_0_in = PE_wrapper295_U0_fifo_w_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] w_IO_L2_in148_U0_fifo_w_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    w_IO_L2_in148_U0_fifo_w_out_V_V_din_pass_0_q0 <= w_IO_L2_in148_U0_fifo_w_out_V_V_din_pass_0_out;
  end
  assign w_IO_L2_in148_U0_fifo_w_out_V_V_din_pass_0_in = w_IO_L2_in148_U0_fifo_w_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  w_IO_L2_in148_U0_fifo_w_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    w_IO_L2_in148_U0_fifo_w_out_V_V_write_pass_0_q0 <= w_IO_L2_in148_U0_fifo_w_out_V_V_write_pass_0_out;
  end
  assign w_IO_L2_in148_U0_fifo_w_out_V_V_write_pass_0_in = w_IO_L2_in148_U0_fifo_w_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_13_4_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_13_4_V_V_full_n_pass_0_q0 <= fifo_w_PE_13_4_V_V_full_n_pass_0_out;
  end
  assign fifo_w_PE_13_4_V_V_full_n_pass_0_in = fifo_w_PE_13_4_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg [63:0] cout_drain_IO_L1_out_wrapper417_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper417_U0_fifo_cout_drain_out_V_V_din_pass_0_q0 <= cout_drain_IO_L1_out_wrapper417_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper417_U0_fifo_cout_drain_out_V_V_din_pass_0_in = cout_drain_IO_L1_out_wrapper417_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  cout_drain_IO_L1_out_wrapper417_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper417_U0_fifo_cout_drain_out_V_V_write_pass_0_q0 <= cout_drain_IO_L1_out_wrapper417_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper417_U0_fifo_cout_drain_out_V_V_write_pass_0_in = cout_drain_IO_L1_out_wrapper417_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [31:0] PE_wrapper308_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper308_U0_fifo_cout_drain_out_V_din_pass_0_q0 <= PE_wrapper308_U0_fifo_cout_drain_out_V_din_pass_0_out;
  end
  assign PE_wrapper308_U0_fifo_cout_drain_out_V_din_pass_0_in = PE_wrapper308_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper308_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper308_U0_fifo_cout_drain_out_V_write_pass_0_q0 <= PE_wrapper308_U0_fifo_cout_drain_out_V_write_pass_0_out;
  end
  assign PE_wrapper308_U0_fifo_cout_drain_out_V_write_pass_0_in = PE_wrapper308_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_w_w_IO_L2_in_13_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_w_IO_L2_in_13_V_V_full_n_pass_0_q0 <= fifo_w_w_IO_L2_in_13_V_V_full_n_pass_0_out;
  end
  assign fifo_w_w_IO_L2_in_13_V_V_full_n_pass_0_in = fifo_w_w_IO_L2_in_13_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_12_0_V_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_12_0_V_V_full_n_pass_1_q0 <= fifo_cin_PE_12_0_V_V_full_n_pass_1_out;
  end
  assign fifo_cin_PE_12_0_V_V_full_n_pass_1_in = fifo_cin_PE_12_0_V_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_cout_drain_IO_L1_out_3_14_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_cout_drain_IO_L1_out_3_14_V_V_full_n_pass_0_q0 <= fifo_cout_drain_cout_drain_IO_L1_out_3_14_V_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_cout_drain_IO_L1_out_3_14_V_V_full_n_pass_0_in = fifo_cout_drain_cout_drain_IO_L1_out_3_14_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper297_U0_fifo_cin_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper297_U0_fifo_cin_out_V_V_din_pass_0_q0 <= PE_wrapper297_U0_fifo_cin_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper297_U0_fifo_cin_out_V_V_din_pass_0_in = PE_wrapper297_U0_fifo_cin_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper297_U0_fifo_cin_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper297_U0_fifo_cin_out_V_V_write_pass_0_q0 <= PE_wrapper297_U0_fifo_cin_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper297_U0_fifo_cin_out_V_V_write_pass_0_in = PE_wrapper297_U0_fifo_cin_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_13_1_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_13_1_V_V_full_n_pass_0_q0 <= fifo_w_PE_13_1_V_V_full_n_pass_0_out;
  end
  assign fifo_w_PE_13_1_V_V_full_n_pass_0_in = fifo_w_PE_13_1_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0_q0 <= PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0_in = PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper238_U0_fifo_cin_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper238_U0_fifo_cin_out_V_V_write_pass_0_q0 <= PE_wrapper238_U0_fifo_cin_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper238_U0_fifo_cin_out_V_V_write_pass_0_in = PE_wrapper238_U0_fifo_cin_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0_q0 <= PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0_in = PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper297_U0_fifo_w_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper297_U0_fifo_w_out_V_V_write_pass_0_q0 <= PE_wrapper297_U0_fifo_w_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper297_U0_fifo_w_out_V_V_write_pass_0_in = PE_wrapper297_U0_fifo_w_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [31:0] PE_wrapper294_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper294_U0_fifo_cout_drain_out_V_din_pass_0_q0 <= PE_wrapper294_U0_fifo_cout_drain_out_V_din_pass_0_out;
  end
  assign PE_wrapper294_U0_fifo_cout_drain_out_V_din_pass_0_in = PE_wrapper294_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper294_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper294_U0_fifo_cout_drain_out_V_write_pass_0_q0 <= PE_wrapper294_U0_fifo_cout_drain_out_V_write_pass_0_out;
  end
  assign PE_wrapper294_U0_fifo_cout_drain_out_V_write_pass_0_in = PE_wrapper294_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0_q0 <= PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0_in = PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper310_U0_fifo_cin_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper310_U0_fifo_cin_out_V_V_write_pass_0_q0 <= PE_wrapper310_U0_fifo_cin_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper310_U0_fifo_cin_out_V_V_write_pass_0_in = PE_wrapper310_U0_fifo_cin_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0_q0 <= PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0_in = PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper307_U0_fifo_cin_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper307_U0_fifo_cin_out_V_V_write_pass_0_q0 <= PE_wrapper307_U0_fifo_cin_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper307_U0_fifo_cin_out_V_V_write_pass_0_in = PE_wrapper307_U0_fifo_cin_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_7_4_V_V_full_n_pass_2_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_7_4_V_V_full_n_pass_2_q0 <= fifo_w_PE_7_4_V_V_full_n_pass_2_out;
  end
  assign fifo_w_PE_7_4_V_V_full_n_pass_2_in = fifo_w_PE_7_4_V_V_full_n_pass_2_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_12_1_V_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_12_1_V_V_full_n_pass_1_q0 <= fifo_cin_PE_12_1_V_V_full_n_pass_1_out;
  end
  assign fifo_cin_PE_12_1_V_V_full_n_pass_1_in = fifo_cin_PE_12_1_V_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg [31:0] PE_wrapper295_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper295_U0_fifo_cout_drain_out_V_din_pass_0_q0 <= PE_wrapper295_U0_fifo_cout_drain_out_V_din_pass_0_out;
  end
  assign PE_wrapper295_U0_fifo_cout_drain_out_V_din_pass_0_in = PE_wrapper295_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper295_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper295_U0_fifo_cout_drain_out_V_write_pass_0_q0 <= PE_wrapper295_U0_fifo_cout_drain_out_V_write_pass_0_out;
  end
  assign PE_wrapper295_U0_fifo_cout_drain_out_V_write_pass_0_in = PE_wrapper295_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper294_U0_fifo_cin_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper294_U0_fifo_cin_out_V_V_din_pass_0_q0 <= PE_wrapper294_U0_fifo_cin_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper294_U0_fifo_cin_out_V_V_din_pass_0_in = PE_wrapper294_U0_fifo_cin_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper294_U0_fifo_cin_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper294_U0_fifo_cin_out_V_V_write_pass_0_q0 <= PE_wrapper294_U0_fifo_cin_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper294_U0_fifo_cin_out_V_V_write_pass_0_in = PE_wrapper294_U0_fifo_cin_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_12_0_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_12_0_V_V_full_n_pass_0_q0 <= fifo_w_PE_12_0_V_V_full_n_pass_0_out;
  end
  assign fifo_w_PE_12_0_V_V_full_n_pass_0_in = fifo_w_PE_12_0_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_cout_drain_IO_L1_out_4_9_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_cout_drain_IO_L1_out_4_9_V_V_full_n_pass_0_q0 <= fifo_cout_drain_cout_drain_IO_L1_out_4_9_V_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_cout_drain_IO_L1_out_4_9_V_V_full_n_pass_0_in = fifo_cout_drain_cout_drain_IO_L1_out_4_9_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg [31:0] PE_wrapper297_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper297_U0_fifo_cout_drain_out_V_din_pass_0_q0 <= PE_wrapper297_U0_fifo_cout_drain_out_V_din_pass_0_out;
  end
  assign PE_wrapper297_U0_fifo_cout_drain_out_V_din_pass_0_in = PE_wrapper297_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper297_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper297_U0_fifo_cout_drain_out_V_write_pass_0_q0 <= PE_wrapper297_U0_fifo_cout_drain_out_V_write_pass_0_out;
  end
  assign PE_wrapper297_U0_fifo_cout_drain_out_V_write_pass_0_in = PE_wrapper297_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper308_U0_fifo_cin_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper308_U0_fifo_cin_out_V_V_din_pass_0_q0 <= PE_wrapper308_U0_fifo_cin_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper308_U0_fifo_cin_out_V_V_din_pass_0_in = PE_wrapper308_U0_fifo_cin_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper308_U0_fifo_cin_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper308_U0_fifo_cin_out_V_V_write_pass_0_q0 <= PE_wrapper308_U0_fifo_cin_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper308_U0_fifo_cin_out_V_V_write_pass_0_in = PE_wrapper308_U0_fifo_cin_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_cout_drain_IO_L1_out_1_14_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_cout_drain_IO_L1_out_1_14_V_V_full_n_pass_0_q0 <= fifo_cout_drain_cout_drain_IO_L1_out_1_14_V_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_cout_drain_IO_L1_out_1_14_V_V_full_n_pass_0_in = fifo_cout_drain_cout_drain_IO_L1_out_1_14_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper308_U0_fifo_w_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper308_U0_fifo_w_out_V_V_din_pass_0_q0 <= PE_wrapper308_U0_fifo_w_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper308_U0_fifo_w_out_V_V_din_pass_0_in = PE_wrapper308_U0_fifo_w_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper308_U0_fifo_w_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper308_U0_fifo_w_out_V_V_write_pass_0_q0 <= PE_wrapper308_U0_fifo_w_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper308_U0_fifo_w_out_V_V_write_pass_0_in = PE_wrapper308_U0_fifo_w_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_13_2_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_13_2_V_V_full_n_pass_0_q0 <= fifo_cin_PE_13_2_V_V_full_n_pass_0_out;
  end
  assign fifo_cin_PE_13_2_V_V_full_n_pass_0_in = fifo_cin_PE_13_2_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_12_3_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_12_3_V_V_full_n_pass_0_q0 <= fifo_w_PE_12_3_V_V_full_n_pass_0_out;
  end
  assign fifo_w_PE_12_3_V_V_full_n_pass_0_in = fifo_w_PE_12_3_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_7_4_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_7_4_V_V_full_n_pass_0_q0 <= fifo_cin_PE_7_4_V_V_full_n_pass_0_out;
  end
  assign fifo_cin_PE_7_4_V_V_full_n_pass_0_in = fifo_cin_PE_7_4_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] w_IO_L2_in148_U0_fifo_w_local_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    w_IO_L2_in148_U0_fifo_w_local_out_V_V_din_pass_0_q0 <= w_IO_L2_in148_U0_fifo_w_local_out_V_V_din_pass_0_out;
  end
  assign w_IO_L2_in148_U0_fifo_w_local_out_V_V_din_pass_0_in = w_IO_L2_in148_U0_fifo_w_local_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  w_IO_L2_in148_U0_fifo_w_local_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    w_IO_L2_in148_U0_fifo_w_local_out_V_V_write_pass_0_q0 <= w_IO_L2_in148_U0_fifo_w_local_out_V_V_write_pass_0_out;
  end
  assign w_IO_L2_in148_U0_fifo_w_local_out_V_V_write_pass_0_in = w_IO_L2_in148_U0_fifo_w_local_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0_q0 <= PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0_in = PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper238_U0_fifo_w_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper238_U0_fifo_w_out_V_V_write_pass_0_q0 <= PE_wrapper238_U0_fifo_w_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper238_U0_fifo_w_out_V_V_write_pass_0_in = PE_wrapper238_U0_fifo_w_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_12_3_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_12_3_V_V_full_n_pass_0_q0 <= fifo_cin_PE_12_3_V_V_full_n_pass_0_out;
  end
  assign fifo_cin_PE_12_3_V_V_full_n_pass_0_in = fifo_cin_PE_12_3_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_PE_13_3_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_PE_13_3_V_full_n_pass_0_q0 <= fifo_cout_drain_PE_13_3_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_PE_13_3_V_full_n_pass_0_in = fifo_cout_drain_PE_13_3_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  ap_done_Boundary_X0Y6_To_X2Y6_q0;
  always @ (posedge ap_clk) begin
    ap_done_Boundary_X0Y6_To_X2Y6_q0 <= ap_done_Boundary_X0Y6_To_X2Y6_out;
  end
  assign ap_done_Boundary_X0Y6_To_X2Y6_in = ap_done_Boundary_X0Y6_To_X2Y6_q0;
  (* dont_touch = "yes" *) reg  ap_start_Boundary_X0Y8_To_X2Y8_q0;
  always @ (posedge ap_clk) begin
    ap_start_Boundary_X0Y8_To_X2Y8_q0 <= ap_start_Boundary_X0Y8_To_X2Y8_out;
  end
  assign ap_start_Boundary_X0Y8_To_X2Y8_in = ap_start_Boundary_X0Y8_To_X2Y8_q0;
  (* dont_touch = "yes" *) reg  ap_rst_n_Boundary_X0Y8_To_X2Y8_q0;
  always @ (posedge ap_clk) begin
    ap_rst_n_Boundary_X0Y8_To_X2Y8_q0 <= ap_rst_n_Boundary_X0Y8_To_X2Y8_out;
  end
  assign ap_rst_n_Boundary_X0Y8_To_X2Y8_in = ap_rst_n_Boundary_X0Y8_To_X2Y8_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper309_U0_fifo_cin_out_V_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper309_U0_fifo_cin_out_V_V_din_pass_1_q0 <= PE_wrapper309_U0_fifo_cin_out_V_V_din_pass_1_out;
  end
  assign PE_wrapper309_U0_fifo_cin_out_V_V_din_pass_1_in = PE_wrapper309_U0_fifo_cin_out_V_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_14_3_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_14_3_V_V_full_n_pass_0_q0 <= fifo_cin_PE_14_3_V_V_full_n_pass_0_out;
  end
  assign fifo_cin_PE_14_3_V_V_full_n_pass_0_in = fifo_cin_PE_14_3_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper309_U0_fifo_cin_out_V_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper309_U0_fifo_cin_out_V_V_write_pass_1_q0 <= PE_wrapper309_U0_fifo_cin_out_V_V_write_pass_1_out;
  end
  assign PE_wrapper309_U0_fifo_cin_out_V_V_write_pass_1_in = PE_wrapper309_U0_fifo_cin_out_V_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper214_U0_fifo_cin_out_V_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper214_U0_fifo_cin_out_V_V_din_pass_1_q0 <= PE_wrapper214_U0_fifo_cin_out_V_V_din_pass_1_out;
  end
  assign PE_wrapper214_U0_fifo_cin_out_V_V_din_pass_1_in = PE_wrapper214_U0_fifo_cin_out_V_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_6_4_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_6_4_V_V_full_n_pass_0_q0 <= fifo_cin_PE_6_4_V_V_full_n_pass_0_out;
  end
  assign fifo_cin_PE_6_4_V_V_full_n_pass_0_in = fifo_cin_PE_6_4_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper214_U0_fifo_cin_out_V_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper214_U0_fifo_cin_out_V_V_write_pass_1_q0 <= PE_wrapper214_U0_fifo_cin_out_V_V_write_pass_1_out;
  end
  assign PE_wrapper214_U0_fifo_cin_out_V_V_write_pass_1_in = PE_wrapper214_U0_fifo_cin_out_V_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [63:0] cout_drain_IO_L1_out_wrapper418_U0_fifo_cout_drain_out_V_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper418_U0_fifo_cout_drain_out_V_V_din_pass_1_q0 <= cout_drain_IO_L1_out_wrapper418_U0_fifo_cout_drain_out_V_V_din_pass_1_out;
  end
  assign cout_drain_IO_L1_out_wrapper418_U0_fifo_cout_drain_out_V_V_din_pass_1_in = cout_drain_IO_L1_out_wrapper418_U0_fifo_cout_drain_out_V_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_cout_drain_IO_L1_out_3_12_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_cout_drain_IO_L1_out_3_12_V_V_full_n_pass_0_q0 <= fifo_cout_drain_cout_drain_IO_L1_out_3_12_V_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_cout_drain_IO_L1_out_3_12_V_V_full_n_pass_0_in = fifo_cout_drain_cout_drain_IO_L1_out_3_12_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  cout_drain_IO_L1_out_wrapper418_U0_fifo_cout_drain_out_V_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper418_U0_fifo_cout_drain_out_V_V_write_pass_1_q0 <= cout_drain_IO_L1_out_wrapper418_U0_fifo_cout_drain_out_V_V_write_pass_1_out;
  end
  assign cout_drain_IO_L1_out_wrapper418_U0_fifo_cout_drain_out_V_V_write_pass_1_in = cout_drain_IO_L1_out_wrapper418_U0_fifo_cout_drain_out_V_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper225_U0_fifo_w_out_V_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper225_U0_fifo_w_out_V_V_din_pass_1_q0 <= PE_wrapper225_U0_fifo_w_out_V_V_din_pass_1_out;
  end
  assign PE_wrapper225_U0_fifo_w_out_V_V_din_pass_1_in = PE_wrapper225_U0_fifo_w_out_V_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_6_4_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_6_4_V_V_full_n_pass_0_q0 <= fifo_w_PE_6_4_V_V_full_n_pass_0_out;
  end
  assign fifo_w_PE_6_4_V_V_full_n_pass_0_in = fifo_w_PE_6_4_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper225_U0_fifo_w_out_V_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper225_U0_fifo_w_out_V_V_write_pass_1_q0 <= PE_wrapper225_U0_fifo_w_out_V_V_write_pass_1_out;
  end
  assign PE_wrapper225_U0_fifo_w_out_V_V_write_pass_1_in = PE_wrapper225_U0_fifo_w_out_V_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper285_U0_fifo_w_out_V_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper285_U0_fifo_w_out_V_V_din_pass_1_q0 <= PE_wrapper285_U0_fifo_w_out_V_V_din_pass_1_out;
  end
  assign PE_wrapper285_U0_fifo_w_out_V_V_din_pass_1_in = PE_wrapper285_U0_fifo_w_out_V_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_11_4_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_11_4_V_V_full_n_pass_0_q0 <= fifo_w_PE_11_4_V_V_full_n_pass_0_out;
  end
  assign fifo_w_PE_11_4_V_V_full_n_pass_0_in = fifo_w_PE_11_4_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper285_U0_fifo_w_out_V_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper285_U0_fifo_w_out_V_V_write_pass_1_q0 <= PE_wrapper285_U0_fifo_w_out_V_V_write_pass_1_out;
  end
  assign PE_wrapper285_U0_fifo_w_out_V_V_write_pass_1_in = PE_wrapper285_U0_fifo_w_out_V_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper306_U0_fifo_cin_out_V_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper306_U0_fifo_cin_out_V_V_din_pass_1_q0 <= PE_wrapper306_U0_fifo_cin_out_V_V_din_pass_1_out;
  end
  assign PE_wrapper306_U0_fifo_cin_out_V_V_din_pass_1_in = PE_wrapper306_U0_fifo_cin_out_V_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_14_0_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_14_0_V_V_full_n_pass_0_q0 <= fifo_cin_PE_14_0_V_V_full_n_pass_0_out;
  end
  assign fifo_cin_PE_14_0_V_V_full_n_pass_0_in = fifo_cin_PE_14_0_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper306_U0_fifo_cin_out_V_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper306_U0_fifo_cin_out_V_V_write_pass_1_q0 <= PE_wrapper306_U0_fifo_cin_out_V_V_write_pass_1_out;
  end
  assign PE_wrapper306_U0_fifo_cin_out_V_V_write_pass_1_in = PE_wrapper306_U0_fifo_cin_out_V_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [31:0] PE_wrapper285_U0_fifo_cout_drain_out_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper285_U0_fifo_cout_drain_out_V_din_pass_1_q0 <= PE_wrapper285_U0_fifo_cout_drain_out_V_din_pass_1_out;
  end
  assign PE_wrapper285_U0_fifo_cout_drain_out_V_din_pass_1_in = PE_wrapper285_U0_fifo_cout_drain_out_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_PE_11_3_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_PE_11_3_V_full_n_pass_0_q0 <= fifo_cout_drain_PE_11_3_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_PE_11_3_V_full_n_pass_0_in = fifo_cout_drain_PE_11_3_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper285_U0_fifo_cout_drain_out_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper285_U0_fifo_cout_drain_out_V_write_pass_1_q0 <= PE_wrapper285_U0_fifo_cout_drain_out_V_write_pass_1_out;
  end
  assign PE_wrapper285_U0_fifo_cout_drain_out_V_write_pass_1_in = PE_wrapper285_U0_fifo_cout_drain_out_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper262_U0_fifo_cin_out_V_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper262_U0_fifo_cin_out_V_V_din_pass_1_q0 <= PE_wrapper262_U0_fifo_cin_out_V_V_din_pass_1_out;
  end
  assign PE_wrapper262_U0_fifo_cin_out_V_V_din_pass_1_in = PE_wrapper262_U0_fifo_cin_out_V_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_10_4_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_10_4_V_V_full_n_pass_0_q0 <= fifo_cin_PE_10_4_V_V_full_n_pass_0_out;
  end
  assign fifo_cin_PE_10_4_V_V_full_n_pass_0_in = fifo_cin_PE_10_4_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper262_U0_fifo_cin_out_V_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper262_U0_fifo_cin_out_V_V_write_pass_1_q0 <= PE_wrapper262_U0_fifo_cin_out_V_V_write_pass_1_out;
  end
  assign PE_wrapper262_U0_fifo_cin_out_V_V_write_pass_1_in = PE_wrapper262_U0_fifo_cin_out_V_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [31:0] PE_wrapper296_U0_fifo_cout_drain_out_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper296_U0_fifo_cout_drain_out_V_din_pass_1_q0 <= PE_wrapper296_U0_fifo_cout_drain_out_V_din_pass_1_out;
  end
  assign PE_wrapper296_U0_fifo_cout_drain_out_V_din_pass_1_in = PE_wrapper296_U0_fifo_cout_drain_out_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_PE_12_2_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_PE_12_2_V_full_n_pass_0_q0 <= fifo_cout_drain_PE_12_2_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_PE_12_2_V_full_n_pass_0_in = fifo_cout_drain_PE_12_2_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper296_U0_fifo_cout_drain_out_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper296_U0_fifo_cout_drain_out_V_write_pass_1_q0 <= PE_wrapper296_U0_fifo_cout_drain_out_V_write_pass_1_out;
  end
  assign PE_wrapper296_U0_fifo_cout_drain_out_V_write_pass_1_in = PE_wrapper296_U0_fifo_cout_drain_out_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [63:0] cout_drain_IO_L1_out_wrapper440_U0_fifo_cout_drain_out_V_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper440_U0_fifo_cout_drain_out_V_V_din_pass_1_q0 <= cout_drain_IO_L1_out_wrapper440_U0_fifo_cout_drain_out_V_V_din_pass_1_out;
  end
  assign cout_drain_IO_L1_out_wrapper440_U0_fifo_cout_drain_out_V_V_din_pass_1_in = cout_drain_IO_L1_out_wrapper440_U0_fifo_cout_drain_out_V_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_cout_drain_IO_L1_out_4_6_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_cout_drain_IO_L1_out_4_6_V_V_full_n_pass_0_q0 <= fifo_cout_drain_cout_drain_IO_L1_out_4_6_V_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_cout_drain_IO_L1_out_4_6_V_V_full_n_pass_0_in = fifo_cout_drain_cout_drain_IO_L1_out_4_6_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  cout_drain_IO_L1_out_wrapper440_U0_fifo_cout_drain_out_V_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper440_U0_fifo_cout_drain_out_V_V_write_pass_1_q0 <= cout_drain_IO_L1_out_wrapper440_U0_fifo_cout_drain_out_V_V_write_pass_1_out;
  end
  assign cout_drain_IO_L1_out_wrapper440_U0_fifo_cout_drain_out_V_V_write_pass_1_in = cout_drain_IO_L1_out_wrapper440_U0_fifo_cout_drain_out_V_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_PE_14_2_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_PE_14_2_V_full_n_pass_0_q0 <= fifo_cout_drain_PE_14_2_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_PE_14_2_V_full_n_pass_0_in = fifo_cout_drain_PE_14_2_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg [63:0] cout_drain_IO_L1_out_wrapper433_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper433_U0_fifo_cout_drain_out_V_V_din_pass_0_q0 <= cout_drain_IO_L1_out_wrapper433_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper433_U0_fifo_cout_drain_out_V_V_din_pass_0_in = cout_drain_IO_L1_out_wrapper433_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  cout_drain_IO_L1_out_wrapper433_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper433_U0_fifo_cout_drain_out_V_V_write_pass_0_q0 <= cout_drain_IO_L1_out_wrapper433_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper433_U0_fifo_cout_drain_out_V_V_write_pass_0_in = cout_drain_IO_L1_out_wrapper433_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_15_4_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_15_4_V_V_full_n_pass_0_q0 <= fifo_w_PE_15_4_V_V_full_n_pass_0_out;
  end
  assign fifo_w_PE_15_4_V_V_full_n_pass_0_in = fifo_w_PE_15_4_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_w_w_IO_L2_in_15_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_w_IO_L2_in_15_V_V_full_n_pass_0_q0 <= fifo_w_w_IO_L2_in_15_V_V_full_n_pass_0_out;
  end
  assign fifo_w_w_IO_L2_in_15_V_V_full_n_pass_0_in = fifo_w_w_IO_L2_in_15_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper250_U0_fifo_cin_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper250_U0_fifo_cin_out_V_V_din_pass_0_q0 <= PE_wrapper250_U0_fifo_cin_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper250_U0_fifo_cin_out_V_V_din_pass_0_in = PE_wrapper250_U0_fifo_cin_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper250_U0_fifo_cin_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper250_U0_fifo_cin_out_V_V_write_pass_0_q0 <= PE_wrapper250_U0_fifo_cin_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper250_U0_fifo_cin_out_V_V_write_pass_0_in = PE_wrapper250_U0_fifo_cin_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [31:0] PE_wrapper250_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper250_U0_fifo_cout_drain_out_V_din_pass_0_q0 <= PE_wrapper250_U0_fifo_cout_drain_out_V_din_pass_0_out;
  end
  assign PE_wrapper250_U0_fifo_cout_drain_out_V_din_pass_0_in = PE_wrapper250_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper250_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper250_U0_fifo_cout_drain_out_V_write_pass_0_q0 <= PE_wrapper250_U0_fifo_cout_drain_out_V_write_pass_0_out;
  end
  assign PE_wrapper250_U0_fifo_cout_drain_out_V_write_pass_0_in = PE_wrapper250_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper298_U0_fifo_cin_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper298_U0_fifo_cin_out_V_V_din_pass_0_q0 <= PE_wrapper298_U0_fifo_cin_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper298_U0_fifo_cin_out_V_V_din_pass_0_in = PE_wrapper298_U0_fifo_cin_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper298_U0_fifo_cin_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper298_U0_fifo_cin_out_V_V_write_pass_0_q0 <= PE_wrapper298_U0_fifo_cin_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper298_U0_fifo_cin_out_V_V_write_pass_0_in = PE_wrapper298_U0_fifo_cin_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_cout_drain_IO_L1_out_4_14_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_cout_drain_IO_L1_out_4_14_V_V_full_n_pass_0_q0 <= fifo_cout_drain_cout_drain_IO_L1_out_4_14_V_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_cout_drain_IO_L1_out_4_14_V_V_full_n_pass_0_in = fifo_cout_drain_cout_drain_IO_L1_out_4_14_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_14_1_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_14_1_V_V_full_n_pass_0_q0 <= fifo_w_PE_14_1_V_V_full_n_pass_0_out;
  end
  assign fifo_w_PE_14_1_V_V_full_n_pass_0_in = fifo_w_PE_14_1_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_PE_13_0_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_PE_13_0_V_full_n_pass_0_q0 <= fifo_cout_drain_PE_13_0_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_PE_13_0_V_full_n_pass_0_in = fifo_cout_drain_PE_13_0_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_PE_13_4_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_PE_13_4_V_full_n_pass_1_q0 <= fifo_cout_drain_PE_13_4_V_full_n_pass_1_out;
  end
  assign fifo_cout_drain_PE_13_4_V_full_n_pass_1_in = fifo_cout_drain_PE_13_4_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_12_4_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_12_4_V_V_full_n_pass_0_q0 <= fifo_cin_PE_12_4_V_V_full_n_pass_0_out;
  end
  assign fifo_cin_PE_12_4_V_V_full_n_pass_0_in = fifo_cin_PE_12_4_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper331_U0_fifo_w_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper331_U0_fifo_w_out_V_V_din_pass_0_q0 <= PE_wrapper331_U0_fifo_w_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper331_U0_fifo_w_out_V_V_din_pass_0_in = PE_wrapper331_U0_fifo_w_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper331_U0_fifo_w_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper331_U0_fifo_w_out_V_V_write_pass_0_q0 <= PE_wrapper331_U0_fifo_w_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper331_U0_fifo_w_out_V_V_write_pass_0_in = PE_wrapper331_U0_fifo_w_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_PE_13_2_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_PE_13_2_V_full_n_pass_1_q0 <= fifo_cout_drain_PE_13_2_V_full_n_pass_1_out;
  end
  assign fifo_cout_drain_PE_13_2_V_full_n_pass_1_in = fifo_cout_drain_PE_13_2_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_15_1_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_15_1_V_V_full_n_pass_0_q0 <= fifo_w_PE_15_1_V_V_full_n_pass_0_out;
  end
  assign fifo_w_PE_15_1_V_V_full_n_pass_0_in = fifo_w_PE_15_1_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_16_0_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_16_0_V_V_full_n_pass_0_q0 <= fifo_cin_PE_16_0_V_V_full_n_pass_0_out;
  end
  assign fifo_cin_PE_16_0_V_V_full_n_pass_0_in = fifo_cin_PE_16_0_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_cout_drain_IO_L1_out_3_11_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_cout_drain_IO_L1_out_3_11_V_V_full_n_pass_0_q0 <= fifo_cout_drain_cout_drain_IO_L1_out_3_11_V_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_cout_drain_IO_L1_out_3_11_V_V_full_n_pass_0_in = fifo_cout_drain_cout_drain_IO_L1_out_3_11_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] w_IO_L2_in_boundary_U0_fifo_w_local_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    w_IO_L2_in_boundary_U0_fifo_w_local_out_V_V_din_pass_0_q0 <= w_IO_L2_in_boundary_U0_fifo_w_local_out_V_V_din_pass_0_out;
  end
  assign w_IO_L2_in_boundary_U0_fifo_w_local_out_V_V_din_pass_0_in = w_IO_L2_in_boundary_U0_fifo_w_local_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  w_IO_L2_in_boundary_U0_fifo_w_local_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    w_IO_L2_in_boundary_U0_fifo_w_local_out_V_V_write_pass_0_q0 <= w_IO_L2_in_boundary_U0_fifo_w_local_out_V_V_write_pass_0_out;
  end
  assign w_IO_L2_in_boundary_U0_fifo_w_local_out_V_V_write_pass_0_in = w_IO_L2_in_boundary_U0_fifo_w_local_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_PE_15_3_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_PE_15_3_V_full_n_pass_0_q0 <= fifo_cout_drain_PE_15_3_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_PE_15_3_V_full_n_pass_0_in = fifo_cout_drain_PE_15_3_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_8_4_V_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_8_4_V_V_full_n_pass_1_q0 <= fifo_cin_PE_8_4_V_V_full_n_pass_1_out;
  end
  assign fifo_cin_PE_8_4_V_V_full_n_pass_1_in = fifo_cin_PE_8_4_V_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_12_4_V_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_12_4_V_V_full_n_pass_1_q0 <= fifo_w_PE_12_4_V_V_full_n_pass_1_out;
  end
  assign fifo_w_PE_12_4_V_V_full_n_pass_1_in = fifo_w_PE_12_4_V_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper273_U0_fifo_w_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper273_U0_fifo_w_out_V_V_din_pass_0_q0 <= PE_wrapper273_U0_fifo_w_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper273_U0_fifo_w_out_V_V_din_pass_0_in = PE_wrapper273_U0_fifo_w_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper273_U0_fifo_w_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper273_U0_fifo_w_out_V_V_write_pass_0_q0 <= PE_wrapper273_U0_fifo_w_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper273_U0_fifo_w_out_V_V_write_pass_0_in = PE_wrapper273_U0_fifo_w_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_14_4_V_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_14_4_V_V_full_n_pass_1_q0 <= fifo_cin_PE_14_4_V_V_full_n_pass_1_out;
  end
  assign fifo_cin_PE_14_4_V_V_full_n_pass_1_in = fifo_cin_PE_14_4_V_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg [63:0] cout_drain_IO_L1_out_boundary_wrapper383_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_boundary_wrapper383_U0_fifo_cout_drain_out_V_V_din_pass_0_q0 <= cout_drain_IO_L1_out_boundary_wrapper383_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  end
  assign cout_drain_IO_L1_out_boundary_wrapper383_U0_fifo_cout_drain_out_V_V_din_pass_0_in = cout_drain_IO_L1_out_boundary_wrapper383_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  cout_drain_IO_L1_out_boundary_wrapper383_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_boundary_wrapper383_U0_fifo_cout_drain_out_V_V_write_pass_0_q0 <= cout_drain_IO_L1_out_boundary_wrapper383_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  end
  assign cout_drain_IO_L1_out_boundary_wrapper383_U0_fifo_cout_drain_out_V_V_write_pass_0_in = cout_drain_IO_L1_out_boundary_wrapper383_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_14_1_V_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_14_1_V_V_full_n_pass_1_q0 <= fifo_cin_PE_14_1_V_V_full_n_pass_1_out;
  end
  assign fifo_cin_PE_14_1_V_V_full_n_pass_1_in = fifo_cin_PE_14_1_V_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_PE_15_0_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_PE_15_0_V_full_n_pass_0_q0 <= fifo_cout_drain_PE_15_0_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_PE_15_0_V_full_n_pass_0_in = fifo_cout_drain_PE_15_0_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0_q0 <= PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0_in = PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper250_U0_fifo_w_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper250_U0_fifo_w_out_V_V_write_pass_0_q0 <= PE_wrapper250_U0_fifo_w_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper250_U0_fifo_w_out_V_V_write_pass_0_in = PE_wrapper250_U0_fifo_w_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper273_U0_fifo_cin_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper273_U0_fifo_cin_out_V_V_din_pass_0_q0 <= PE_wrapper273_U0_fifo_cin_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper273_U0_fifo_cin_out_V_V_din_pass_0_in = PE_wrapper273_U0_fifo_cin_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper273_U0_fifo_cin_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper273_U0_fifo_cin_out_V_V_write_pass_0_q0 <= PE_wrapper273_U0_fifo_cin_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper273_U0_fifo_cin_out_V_V_write_pass_0_in = PE_wrapper273_U0_fifo_cin_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [63:0] cout_drain_IO_L1_out_wrapper369_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper369_U0_fifo_cout_drain_out_V_V_din_pass_0_q0 <= cout_drain_IO_L1_out_wrapper369_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper369_U0_fifo_cout_drain_out_V_V_din_pass_0_in = cout_drain_IO_L1_out_wrapper369_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  cout_drain_IO_L1_out_wrapper369_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper369_U0_fifo_cout_drain_out_V_V_write_pass_0_q0 <= cout_drain_IO_L1_out_wrapper369_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper369_U0_fifo_cout_drain_out_V_V_write_pass_0_in = cout_drain_IO_L1_out_wrapper369_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper319_U0_fifo_w_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper319_U0_fifo_w_out_V_V_din_pass_0_q0 <= PE_wrapper319_U0_fifo_w_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper319_U0_fifo_w_out_V_V_din_pass_0_in = PE_wrapper319_U0_fifo_w_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper319_U0_fifo_w_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper319_U0_fifo_w_out_V_V_write_pass_0_q0 <= PE_wrapper319_U0_fifo_w_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper319_U0_fifo_w_out_V_V_write_pass_0_in = PE_wrapper319_U0_fifo_w_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_8_4_V_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_8_4_V_V_full_n_pass_1_q0 <= fifo_w_PE_8_4_V_V_full_n_pass_1_out;
  end
  assign fifo_w_PE_8_4_V_V_full_n_pass_1_in = fifo_w_PE_8_4_V_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg [31:0] PE_wrapper319_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper319_U0_fifo_cout_drain_out_V_din_pass_0_q0 <= PE_wrapper319_U0_fifo_cout_drain_out_V_din_pass_0_out;
  end
  assign PE_wrapper319_U0_fifo_cout_drain_out_V_din_pass_0_in = PE_wrapper319_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper319_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper319_U0_fifo_cout_drain_out_V_write_pass_0_q0 <= PE_wrapper319_U0_fifo_cout_drain_out_V_write_pass_0_out;
  end
  assign PE_wrapper319_U0_fifo_cout_drain_out_V_write_pass_0_in = PE_wrapper319_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper298_U0_fifo_w_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper298_U0_fifo_w_out_V_V_din_pass_0_q0 <= PE_wrapper298_U0_fifo_w_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper298_U0_fifo_w_out_V_V_din_pass_0_in = PE_wrapper298_U0_fifo_w_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper298_U0_fifo_w_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper298_U0_fifo_w_out_V_V_write_pass_0_q0 <= PE_wrapper298_U0_fifo_w_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper298_U0_fifo_w_out_V_V_write_pass_0_in = PE_wrapper298_U0_fifo_w_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [31:0] PE_wrapper334_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper334_U0_fifo_cout_drain_out_V_din_pass_0_q0 <= PE_wrapper334_U0_fifo_cout_drain_out_V_din_pass_0_out;
  end
  assign PE_wrapper334_U0_fifo_cout_drain_out_V_din_pass_0_in = PE_wrapper334_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper334_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper334_U0_fifo_cout_drain_out_V_write_pass_0_q0 <= PE_wrapper334_U0_fifo_cout_drain_out_V_write_pass_0_out;
  end
  assign PE_wrapper334_U0_fifo_cout_drain_out_V_write_pass_0_in = PE_wrapper334_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper322_U0_fifo_w_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper322_U0_fifo_w_out_V_V_din_pass_0_q0 <= PE_wrapper322_U0_fifo_w_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper322_U0_fifo_w_out_V_V_din_pass_0_in = PE_wrapper322_U0_fifo_w_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper322_U0_fifo_w_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper322_U0_fifo_w_out_V_V_write_pass_0_q0 <= PE_wrapper322_U0_fifo_w_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper322_U0_fifo_w_out_V_V_write_pass_0_in = PE_wrapper322_U0_fifo_w_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [63:0] cout_drain_IO_L1_out_boundary_wrapper415_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_boundary_wrapper415_U0_fifo_cout_drain_out_V_V_din_pass_0_q0 <= cout_drain_IO_L1_out_boundary_wrapper415_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  end
  assign cout_drain_IO_L1_out_boundary_wrapper415_U0_fifo_cout_drain_out_V_V_din_pass_0_in = cout_drain_IO_L1_out_boundary_wrapper415_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  cout_drain_IO_L1_out_boundary_wrapper415_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_boundary_wrapper415_U0_fifo_cout_drain_out_V_V_write_pass_0_q0 <= cout_drain_IO_L1_out_boundary_wrapper415_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  end
  assign cout_drain_IO_L1_out_boundary_wrapper415_U0_fifo_cout_drain_out_V_V_write_pass_0_in = cout_drain_IO_L1_out_boundary_wrapper415_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [63:0] cout_drain_IO_L1_out_wrapper420_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper420_U0_fifo_cout_drain_out_V_V_din_pass_0_q0 <= cout_drain_IO_L1_out_wrapper420_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper420_U0_fifo_cout_drain_out_V_V_din_pass_0_in = cout_drain_IO_L1_out_wrapper420_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  cout_drain_IO_L1_out_wrapper420_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper420_U0_fifo_cout_drain_out_V_V_write_pass_0_q0 <= cout_drain_IO_L1_out_wrapper420_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper420_U0_fifo_cout_drain_out_V_V_write_pass_0_in = cout_drain_IO_L1_out_wrapper420_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_PE_14_0_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_PE_14_0_V_full_n_pass_0_q0 <= fifo_cout_drain_PE_14_0_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_PE_14_0_V_full_n_pass_0_in = fifo_cout_drain_PE_14_0_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_14_4_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_14_4_V_V_full_n_pass_0_q0 <= fifo_w_PE_14_4_V_V_full_n_pass_0_out;
  end
  assign fifo_w_PE_14_4_V_V_full_n_pass_0_in = fifo_w_PE_14_4_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg [31:0] PE_wrapper322_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper322_U0_fifo_cout_drain_out_V_din_pass_0_q0 <= PE_wrapper322_U0_fifo_cout_drain_out_V_din_pass_0_out;
  end
  assign PE_wrapper322_U0_fifo_cout_drain_out_V_din_pass_0_in = PE_wrapper322_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper322_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper322_U0_fifo_cout_drain_out_V_write_pass_0_q0 <= PE_wrapper322_U0_fifo_cout_drain_out_V_write_pass_0_out;
  end
  assign PE_wrapper322_U0_fifo_cout_drain_out_V_write_pass_0_in = PE_wrapper322_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper334_U0_fifo_w_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper334_U0_fifo_w_out_V_V_din_pass_0_q0 <= PE_wrapper334_U0_fifo_w_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper334_U0_fifo_w_out_V_V_din_pass_0_in = PE_wrapper334_U0_fifo_w_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper334_U0_fifo_w_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper334_U0_fifo_w_out_V_V_write_pass_0_q0 <= PE_wrapper334_U0_fifo_w_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper334_U0_fifo_w_out_V_V_write_pass_0_in = PE_wrapper334_U0_fifo_w_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_10_3_V_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_10_3_V_V_full_n_pass_1_q0 <= fifo_w_PE_10_3_V_V_full_n_pass_1_out;
  end
  assign fifo_w_PE_10_3_V_V_full_n_pass_1_in = fifo_w_PE_10_3_V_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_10_3_V_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_10_3_V_V_full_n_pass_1_q0 <= fifo_cin_PE_10_3_V_V_full_n_pass_1_out;
  end
  assign fifo_cin_PE_10_3_V_V_full_n_pass_1_in = fifo_cin_PE_10_3_V_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_cout_drain_IO_L1_out_2_15_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_cout_drain_IO_L1_out_2_15_V_V_full_n_pass_0_q0 <= fifo_cout_drain_cout_drain_IO_L1_out_2_15_V_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_cout_drain_IO_L1_out_2_15_V_V_full_n_pass_0_in = fifo_cout_drain_cout_drain_IO_L1_out_2_15_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg [63:0] cout_drain_IO_L1_out_wrapper401_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper401_U0_fifo_cout_drain_out_V_V_din_pass_0_q0 <= cout_drain_IO_L1_out_wrapper401_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper401_U0_fifo_cout_drain_out_V_V_din_pass_0_in = cout_drain_IO_L1_out_wrapper401_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  cout_drain_IO_L1_out_wrapper401_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper401_U0_fifo_cout_drain_out_V_V_write_pass_0_q0 <= cout_drain_IO_L1_out_wrapper401_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper401_U0_fifo_cout_drain_out_V_V_write_pass_0_in = cout_drain_IO_L1_out_wrapper401_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [31:0] PE_wrapper298_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper298_U0_fifo_cout_drain_out_V_din_pass_0_q0 <= PE_wrapper298_U0_fifo_cout_drain_out_V_din_pass_0_out;
  end
  assign PE_wrapper298_U0_fifo_cout_drain_out_V_din_pass_0_in = PE_wrapper298_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper298_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper298_U0_fifo_cout_drain_out_V_write_pass_0_q0 <= PE_wrapper298_U0_fifo_cout_drain_out_V_write_pass_0_out;
  end
  assign PE_wrapper298_U0_fifo_cout_drain_out_V_write_pass_0_in = PE_wrapper298_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  ap_done_Boundary_X2Y4_To_X4Y4_q0;
  always @ (posedge ap_clk) begin
    ap_done_Boundary_X2Y4_To_X4Y4_q0 <= ap_done_Boundary_X2Y4_To_X4Y4_out;
  end
  assign ap_done_Boundary_X2Y4_To_X4Y4_in = ap_done_Boundary_X2Y4_To_X4Y4_q0;
  (* dont_touch = "yes" *) reg  ap_start_Boundary_X2Y6_To_X4Y6_q0;
  always @ (posedge ap_clk) begin
    ap_start_Boundary_X2Y6_To_X4Y6_q0 <= ap_start_Boundary_X2Y6_To_X4Y6_out;
  end
  assign ap_start_Boundary_X2Y6_To_X4Y6_in = ap_start_Boundary_X2Y6_To_X4Y6_q0;
  (* dont_touch = "yes" *) reg  ap_rst_n_Boundary_X2Y6_To_X4Y6_q0;
  always @ (posedge ap_clk) begin
    ap_rst_n_Boundary_X2Y6_To_X4Y6_q0 <= ap_rst_n_Boundary_X2Y6_To_X4Y6_out;
  end
  assign ap_rst_n_Boundary_X2Y6_To_X4Y6_in = ap_rst_n_Boundary_X2Y6_To_X4Y6_q0;
  (* dont_touch = "yes" *) reg [31:0] PE_wrapper310_U0_fifo_cout_drain_out_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper310_U0_fifo_cout_drain_out_V_din_pass_1_q0 <= PE_wrapper310_U0_fifo_cout_drain_out_V_din_pass_1_out;
  end
  assign PE_wrapper310_U0_fifo_cout_drain_out_V_din_pass_1_in = PE_wrapper310_U0_fifo_cout_drain_out_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_PE_13_4_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_PE_13_4_V_full_n_pass_0_q0 <= fifo_cout_drain_PE_13_4_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_PE_13_4_V_full_n_pass_0_in = fifo_cout_drain_PE_13_4_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper310_U0_fifo_cout_drain_out_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper310_U0_fifo_cout_drain_out_V_write_pass_1_q0 <= PE_wrapper310_U0_fifo_cout_drain_out_V_write_pass_1_out;
  end
  assign PE_wrapper310_U0_fifo_cout_drain_out_V_write_pass_1_in = PE_wrapper310_U0_fifo_cout_drain_out_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [31:0] PE_wrapper308_U0_fifo_cout_drain_out_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper308_U0_fifo_cout_drain_out_V_din_pass_1_q0 <= PE_wrapper308_U0_fifo_cout_drain_out_V_din_pass_1_out;
  end
  assign PE_wrapper308_U0_fifo_cout_drain_out_V_din_pass_1_in = PE_wrapper308_U0_fifo_cout_drain_out_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_PE_13_2_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_PE_13_2_V_full_n_pass_0_q0 <= fifo_cout_drain_PE_13_2_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_PE_13_2_V_full_n_pass_0_in = fifo_cout_drain_PE_13_2_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper308_U0_fifo_cout_drain_out_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper308_U0_fifo_cout_drain_out_V_write_pass_1_q0 <= PE_wrapper308_U0_fifo_cout_drain_out_V_write_pass_1_out;
  end
  assign PE_wrapper308_U0_fifo_cout_drain_out_V_write_pass_1_in = PE_wrapper308_U0_fifo_cout_drain_out_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_1_q0 <= PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_1_out;
  end
  assign PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_1_in = PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_8_4_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_8_4_V_V_full_n_pass_0_q0 <= fifo_cin_PE_8_4_V_V_full_n_pass_0_out;
  end
  assign fifo_cin_PE_8_4_V_V_full_n_pass_0_in = fifo_cin_PE_8_4_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper238_U0_fifo_cin_out_V_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper238_U0_fifo_cin_out_V_V_write_pass_1_q0 <= PE_wrapper238_U0_fifo_cin_out_V_V_write_pass_1_out;
  end
  assign PE_wrapper238_U0_fifo_cin_out_V_V_write_pass_1_in = PE_wrapper238_U0_fifo_cin_out_V_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper297_U0_fifo_w_out_V_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper297_U0_fifo_w_out_V_V_din_pass_1_q0 <= PE_wrapper297_U0_fifo_w_out_V_V_din_pass_1_out;
  end
  assign PE_wrapper297_U0_fifo_w_out_V_V_din_pass_1_in = PE_wrapper297_U0_fifo_w_out_V_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_12_4_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_12_4_V_V_full_n_pass_0_q0 <= fifo_w_PE_12_4_V_V_full_n_pass_0_out;
  end
  assign fifo_w_PE_12_4_V_V_full_n_pass_0_in = fifo_w_PE_12_4_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper297_U0_fifo_w_out_V_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper297_U0_fifo_w_out_V_V_write_pass_1_q0 <= PE_wrapper297_U0_fifo_w_out_V_V_write_pass_1_out;
  end
  assign PE_wrapper297_U0_fifo_w_out_V_V_write_pass_1_in = PE_wrapper297_U0_fifo_w_out_V_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_1_q0 <= PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_1_out;
  end
  assign PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_1_in = PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_14_4_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_14_4_V_V_full_n_pass_0_q0 <= fifo_cin_PE_14_4_V_V_full_n_pass_0_out;
  end
  assign fifo_cin_PE_14_4_V_V_full_n_pass_0_in = fifo_cin_PE_14_4_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper310_U0_fifo_cin_out_V_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper310_U0_fifo_cin_out_V_V_write_pass_1_q0 <= PE_wrapper310_U0_fifo_cin_out_V_V_write_pass_1_out;
  end
  assign PE_wrapper310_U0_fifo_cin_out_V_V_write_pass_1_in = PE_wrapper310_U0_fifo_cin_out_V_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_1_q0 <= PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_1_out;
  end
  assign PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_1_in = PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_14_1_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_14_1_V_V_full_n_pass_0_q0 <= fifo_cin_PE_14_1_V_V_full_n_pass_0_out;
  end
  assign fifo_cin_PE_14_1_V_V_full_n_pass_0_in = fifo_cin_PE_14_1_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper307_U0_fifo_cin_out_V_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper307_U0_fifo_cin_out_V_V_write_pass_1_q0 <= PE_wrapper307_U0_fifo_cin_out_V_V_write_pass_1_out;
  end
  assign PE_wrapper307_U0_fifo_cin_out_V_V_write_pass_1_in = PE_wrapper307_U0_fifo_cin_out_V_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper250_U0_fifo_w_out_V_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper250_U0_fifo_w_out_V_V_din_pass_1_q0 <= PE_wrapper250_U0_fifo_w_out_V_V_din_pass_1_out;
  end
  assign PE_wrapper250_U0_fifo_w_out_V_V_din_pass_1_in = PE_wrapper250_U0_fifo_w_out_V_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_8_5_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_8_5_V_V_full_n_pass_0_q0 <= fifo_w_PE_8_5_V_V_full_n_pass_0_out;
  end
  assign fifo_w_PE_8_5_V_V_full_n_pass_0_in = fifo_w_PE_8_5_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper250_U0_fifo_w_out_V_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper250_U0_fifo_w_out_V_V_write_pass_1_q0 <= PE_wrapper250_U0_fifo_w_out_V_V_write_pass_1_out;
  end
  assign PE_wrapper250_U0_fifo_w_out_V_V_write_pass_1_in = PE_wrapper250_U0_fifo_w_out_V_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper238_U0_fifo_w_out_V_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper238_U0_fifo_w_out_V_V_din_pass_1_q0 <= PE_wrapper238_U0_fifo_w_out_V_V_din_pass_1_out;
  end
  assign PE_wrapper238_U0_fifo_w_out_V_V_din_pass_1_in = PE_wrapper238_U0_fifo_w_out_V_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_7_5_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_7_5_V_V_full_n_pass_0_q0 <= fifo_w_PE_7_5_V_V_full_n_pass_0_out;
  end
  assign fifo_w_PE_7_5_V_V_full_n_pass_0_in = fifo_w_PE_7_5_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper238_U0_fifo_w_out_V_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper238_U0_fifo_w_out_V_V_write_pass_1_q0 <= PE_wrapper238_U0_fifo_w_out_V_V_write_pass_1_out;
  end
  assign PE_wrapper238_U0_fifo_w_out_V_V_write_pass_1_in = PE_wrapper238_U0_fifo_w_out_V_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [31:0] PE_wrapper320_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper320_U0_fifo_cout_drain_out_V_din_pass_0_q0 <= PE_wrapper320_U0_fifo_cout_drain_out_V_din_pass_0_out;
  end
  assign PE_wrapper320_U0_fifo_cout_drain_out_V_din_pass_0_in = PE_wrapper320_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper320_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper320_U0_fifo_cout_drain_out_V_write_pass_0_q0 <= PE_wrapper320_U0_fifo_cout_drain_out_V_write_pass_0_out;
  end
  assign PE_wrapper320_U0_fifo_cout_drain_out_V_write_pass_0_in = PE_wrapper320_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_cout_drain_IO_L1_out_4_13_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_cout_drain_IO_L1_out_4_13_V_V_full_n_pass_0_q0 <= fifo_cout_drain_cout_drain_IO_L1_out_4_13_V_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_cout_drain_IO_L1_out_4_13_V_V_full_n_pass_0_in = fifo_cout_drain_cout_drain_IO_L1_out_4_13_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_14_3_V_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_14_3_V_V_full_n_pass_1_q0 <= fifo_cin_PE_14_3_V_V_full_n_pass_1_out;
  end
  assign fifo_cin_PE_14_3_V_V_full_n_pass_1_in = fifo_cin_PE_14_3_V_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg [63:0] cout_drain_IO_L1_out_wrapper402_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper402_U0_fifo_cout_drain_out_V_V_din_pass_0_q0 <= cout_drain_IO_L1_out_wrapper402_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper402_U0_fifo_cout_drain_out_V_V_din_pass_0_in = cout_drain_IO_L1_out_wrapper402_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  cout_drain_IO_L1_out_wrapper402_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper402_U0_fifo_cout_drain_out_V_V_write_pass_0_q0 <= cout_drain_IO_L1_out_wrapper402_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper402_U0_fifo_cout_drain_out_V_V_write_pass_0_in = cout_drain_IO_L1_out_wrapper402_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] w_IO_L2_in149_U0_fifo_w_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    w_IO_L2_in149_U0_fifo_w_out_V_V_din_pass_0_q0 <= w_IO_L2_in149_U0_fifo_w_out_V_V_din_pass_0_out;
  end
  assign w_IO_L2_in149_U0_fifo_w_out_V_V_din_pass_0_in = w_IO_L2_in149_U0_fifo_w_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  w_IO_L2_in149_U0_fifo_w_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    w_IO_L2_in149_U0_fifo_w_out_V_V_write_pass_0_q0 <= w_IO_L2_in149_U0_fifo_w_out_V_V_write_pass_0_out;
  end
  assign w_IO_L2_in149_U0_fifo_w_out_V_V_write_pass_0_in = w_IO_L2_in149_U0_fifo_w_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [31:0] PE_wrapper286_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper286_U0_fifo_cout_drain_out_V_din_pass_0_q0 <= PE_wrapper286_U0_fifo_cout_drain_out_V_din_pass_0_out;
  end
  assign PE_wrapper286_U0_fifo_cout_drain_out_V_din_pass_0_in = PE_wrapper286_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper286_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper286_U0_fifo_cout_drain_out_V_write_pass_0_q0 <= PE_wrapper286_U0_fifo_cout_drain_out_V_write_pass_0_out;
  end
  assign PE_wrapper286_U0_fifo_cout_drain_out_V_write_pass_0_in = PE_wrapper286_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_6_4_V_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_6_4_V_V_full_n_pass_1_q0 <= fifo_cin_PE_6_4_V_V_full_n_pass_1_out;
  end
  assign fifo_cin_PE_6_4_V_V_full_n_pass_1_in = fifo_cin_PE_6_4_V_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg [63:0] cout_drain_IO_L1_out_wrapper432_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper432_U0_fifo_cout_drain_out_V_V_din_pass_0_q0 <= cout_drain_IO_L1_out_wrapper432_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper432_U0_fifo_cout_drain_out_V_V_din_pass_0_in = cout_drain_IO_L1_out_wrapper432_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  cout_drain_IO_L1_out_wrapper432_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper432_U0_fifo_cout_drain_out_V_V_write_pass_0_q0 <= cout_drain_IO_L1_out_wrapper432_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper432_U0_fifo_cout_drain_out_V_V_write_pass_0_in = cout_drain_IO_L1_out_wrapper432_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper318_U0_fifo_w_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper318_U0_fifo_w_out_V_V_din_pass_0_q0 <= PE_wrapper318_U0_fifo_w_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper318_U0_fifo_w_out_V_V_din_pass_0_in = PE_wrapper318_U0_fifo_w_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper318_U0_fifo_w_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper318_U0_fifo_w_out_V_V_write_pass_0_q0 <= PE_wrapper318_U0_fifo_w_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper318_U0_fifo_w_out_V_V_write_pass_0_in = PE_wrapper318_U0_fifo_w_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [31:0] PE_wrapper226_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper226_U0_fifo_cout_drain_out_V_din_pass_0_q0 <= PE_wrapper226_U0_fifo_cout_drain_out_V_din_pass_0_out;
  end
  assign PE_wrapper226_U0_fifo_cout_drain_out_V_din_pass_0_in = PE_wrapper226_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper226_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper226_U0_fifo_cout_drain_out_V_write_pass_0_q0 <= PE_wrapper226_U0_fifo_cout_drain_out_V_write_pass_0_out;
  end
  assign PE_wrapper226_U0_fifo_cout_drain_out_V_write_pass_0_in = PE_wrapper226_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper286_U0_fifo_cin_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper286_U0_fifo_cin_out_V_V_din_pass_0_q0 <= PE_wrapper286_U0_fifo_cin_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper286_U0_fifo_cin_out_V_V_din_pass_0_in = PE_wrapper286_U0_fifo_cin_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper286_U0_fifo_cin_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper286_U0_fifo_cin_out_V_V_write_pass_0_q0 <= PE_wrapper286_U0_fifo_cin_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper286_U0_fifo_cin_out_V_V_write_pass_0_in = PE_wrapper286_U0_fifo_cin_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_w_w_IO_L2_in_14_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_w_IO_L2_in_14_V_V_full_n_pass_0_q0 <= fifo_w_w_IO_L2_in_14_V_V_full_n_pass_0_out;
  end
  assign fifo_w_w_IO_L2_in_14_V_V_full_n_pass_0_in = fifo_w_w_IO_L2_in_14_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper320_U0_fifo_cin_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper320_U0_fifo_cin_out_V_V_din_pass_0_q0 <= PE_wrapper320_U0_fifo_cin_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper320_U0_fifo_cin_out_V_V_din_pass_0_in = PE_wrapper320_U0_fifo_cin_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper320_U0_fifo_cin_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper320_U0_fifo_cin_out_V_V_write_pass_0_q0 <= PE_wrapper320_U0_fifo_cin_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper320_U0_fifo_cin_out_V_V_write_pass_0_in = PE_wrapper320_U0_fifo_cin_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_cout_drain_IO_L1_out_3_12_V_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_cout_drain_IO_L1_out_3_12_V_V_full_n_pass_1_q0 <= fifo_cout_drain_cout_drain_IO_L1_out_3_12_V_V_full_n_pass_1_out;
  end
  assign fifo_cout_drain_cout_drain_IO_L1_out_3_12_V_V_full_n_pass_1_in = fifo_cout_drain_cout_drain_IO_L1_out_3_12_V_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_6_4_V_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_6_4_V_V_full_n_pass_1_q0 <= fifo_w_PE_6_4_V_V_full_n_pass_1_out;
  end
  assign fifo_w_PE_6_4_V_V_full_n_pass_1_in = fifo_w_PE_6_4_V_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg [63:0] cout_drain_IO_L1_out_wrapper416_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper416_U0_fifo_cout_drain_out_V_V_din_pass_0_q0 <= cout_drain_IO_L1_out_wrapper416_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper416_U0_fifo_cout_drain_out_V_V_din_pass_0_in = cout_drain_IO_L1_out_wrapper416_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  cout_drain_IO_L1_out_wrapper416_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper416_U0_fifo_cout_drain_out_V_V_write_pass_0_q0 <= cout_drain_IO_L1_out_wrapper416_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper416_U0_fifo_cout_drain_out_V_V_write_pass_0_in = cout_drain_IO_L1_out_wrapper416_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper330_U0_fifo_cin_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper330_U0_fifo_cin_out_V_V_din_pass_0_q0 <= PE_wrapper330_U0_fifo_cin_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper330_U0_fifo_cin_out_V_V_din_pass_0_in = PE_wrapper330_U0_fifo_cin_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper330_U0_fifo_cin_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper330_U0_fifo_cin_out_V_V_write_pass_0_q0 <= PE_wrapper330_U0_fifo_cin_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper330_U0_fifo_cin_out_V_V_write_pass_0_in = PE_wrapper330_U0_fifo_cin_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper330_U0_fifo_w_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper330_U0_fifo_w_out_V_V_din_pass_0_q0 <= PE_wrapper330_U0_fifo_w_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper330_U0_fifo_w_out_V_V_din_pass_0_in = PE_wrapper330_U0_fifo_w_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper330_U0_fifo_w_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper330_U0_fifo_w_out_V_V_write_pass_0_q0 <= PE_wrapper330_U0_fifo_w_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper330_U0_fifo_w_out_V_V_write_pass_0_in = PE_wrapper330_U0_fifo_w_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_11_4_V_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_11_4_V_V_full_n_pass_1_q0 <= fifo_w_PE_11_4_V_V_full_n_pass_1_out;
  end
  assign fifo_w_PE_11_4_V_V_full_n_pass_1_in = fifo_w_PE_11_4_V_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg [63:0] cout_drain_IO_L1_out_wrapper419_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper419_U0_fifo_cout_drain_out_V_V_din_pass_0_q0 <= cout_drain_IO_L1_out_wrapper419_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper419_U0_fifo_cout_drain_out_V_V_din_pass_0_in = cout_drain_IO_L1_out_wrapper419_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  cout_drain_IO_L1_out_wrapper419_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper419_U0_fifo_cout_drain_out_V_V_write_pass_0_q0 <= cout_drain_IO_L1_out_wrapper419_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper419_U0_fifo_cout_drain_out_V_V_write_pass_0_in = cout_drain_IO_L1_out_wrapper419_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_15_0_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_15_0_V_V_full_n_pass_0_q0 <= fifo_w_PE_15_0_V_V_full_n_pass_0_out;
  end
  assign fifo_w_PE_15_0_V_V_full_n_pass_0_in = fifo_w_PE_15_0_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_10_4_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_10_4_V_V_full_n_pass_0_q0 <= fifo_w_PE_10_4_V_V_full_n_pass_0_out;
  end
  assign fifo_w_PE_10_4_V_V_full_n_pass_0_in = fifo_w_PE_10_4_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper286_U0_fifo_w_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper286_U0_fifo_w_out_V_V_din_pass_0_q0 <= PE_wrapper286_U0_fifo_w_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper286_U0_fifo_w_out_V_V_din_pass_0_in = PE_wrapper286_U0_fifo_w_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper286_U0_fifo_w_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper286_U0_fifo_w_out_V_V_write_pass_0_q0 <= PE_wrapper286_U0_fifo_w_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper286_U0_fifo_w_out_V_V_write_pass_0_in = PE_wrapper286_U0_fifo_w_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_cout_drain_IO_L1_out_1_15_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_cout_drain_IO_L1_out_1_15_V_V_full_n_pass_0_q0 <= fifo_cout_drain_cout_drain_IO_L1_out_1_15_V_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_cout_drain_IO_L1_out_1_15_V_V_full_n_pass_0_in = fifo_cout_drain_cout_drain_IO_L1_out_1_15_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg [31:0] PE_wrapper330_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper330_U0_fifo_cout_drain_out_V_din_pass_0_q0 <= PE_wrapper330_U0_fifo_cout_drain_out_V_din_pass_0_out;
  end
  assign PE_wrapper330_U0_fifo_cout_drain_out_V_din_pass_0_in = PE_wrapper330_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper330_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper330_U0_fifo_cout_drain_out_V_write_pass_0_q0 <= PE_wrapper330_U0_fifo_cout_drain_out_V_write_pass_0_out;
  end
  assign PE_wrapper330_U0_fifo_cout_drain_out_V_write_pass_0_in = PE_wrapper330_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_14_0_V_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_14_0_V_V_full_n_pass_1_q0 <= fifo_cin_PE_14_0_V_V_full_n_pass_1_out;
  end
  assign fifo_cin_PE_14_0_V_V_full_n_pass_1_in = fifo_cin_PE_14_0_V_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper321_U0_fifo_cin_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper321_U0_fifo_cin_out_V_V_din_pass_0_q0 <= PE_wrapper321_U0_fifo_cin_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper321_U0_fifo_cin_out_V_V_din_pass_0_in = PE_wrapper321_U0_fifo_cin_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper321_U0_fifo_cin_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper321_U0_fifo_cin_out_V_V_write_pass_0_q0 <= PE_wrapper321_U0_fifo_cin_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper321_U0_fifo_cin_out_V_V_write_pass_0_in = PE_wrapper321_U0_fifo_cin_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_PE_11_3_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_PE_11_3_V_full_n_pass_1_q0 <= fifo_cout_drain_PE_11_3_V_full_n_pass_1_out;
  end
  assign fifo_cout_drain_PE_11_3_V_full_n_pass_1_in = fifo_cout_drain_PE_11_3_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_14_2_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_14_2_V_V_full_n_pass_0_q0 <= fifo_w_PE_14_2_V_V_full_n_pass_0_out;
  end
  assign fifo_w_PE_14_2_V_V_full_n_pass_0_in = fifo_w_PE_14_2_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper226_U0_fifo_w_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper226_U0_fifo_w_out_V_V_din_pass_0_q0 <= PE_wrapper226_U0_fifo_w_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper226_U0_fifo_w_out_V_V_din_pass_0_in = PE_wrapper226_U0_fifo_w_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper226_U0_fifo_w_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper226_U0_fifo_w_out_V_V_write_pass_0_q0 <= PE_wrapper226_U0_fifo_w_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper226_U0_fifo_w_out_V_V_write_pass_0_in = PE_wrapper226_U0_fifo_w_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_14_2_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_14_2_V_V_full_n_pass_0_q0 <= fifo_cin_PE_14_2_V_V_full_n_pass_0_out;
  end
  assign fifo_cin_PE_14_2_V_V_full_n_pass_0_in = fifo_cin_PE_14_2_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg [63:0] cout_drain_IO_L1_out_wrapper384_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper384_U0_fifo_cout_drain_out_V_V_din_pass_0_q0 <= cout_drain_IO_L1_out_wrapper384_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper384_U0_fifo_cout_drain_out_V_V_din_pass_0_in = cout_drain_IO_L1_out_wrapper384_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  cout_drain_IO_L1_out_wrapper384_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper384_U0_fifo_cout_drain_out_V_V_write_pass_0_q0 <= cout_drain_IO_L1_out_wrapper384_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper384_U0_fifo_cout_drain_out_V_V_write_pass_0_in = cout_drain_IO_L1_out_wrapper384_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_PE_14_1_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_PE_14_1_V_full_n_pass_0_q0 <= fifo_cout_drain_PE_14_1_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_PE_14_1_V_full_n_pass_0_in = fifo_cout_drain_PE_14_1_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_PE_15_4_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_PE_15_4_V_full_n_pass_0_q0 <= fifo_cout_drain_PE_15_4_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_PE_15_4_V_full_n_pass_0_in = fifo_cout_drain_PE_15_4_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_cout_drain_IO_L1_out_3_15_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_cout_drain_IO_L1_out_3_15_V_V_full_n_pass_0_q0 <= fifo_cout_drain_cout_drain_IO_L1_out_3_15_V_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_cout_drain_IO_L1_out_3_15_V_V_full_n_pass_0_in = fifo_cout_drain_cout_drain_IO_L1_out_3_15_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper274_U0_fifo_w_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper274_U0_fifo_w_out_V_V_din_pass_0_q0 <= PE_wrapper274_U0_fifo_w_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper274_U0_fifo_w_out_V_V_din_pass_0_in = PE_wrapper274_U0_fifo_w_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper274_U0_fifo_w_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper274_U0_fifo_w_out_V_V_write_pass_0_q0 <= PE_wrapper274_U0_fifo_w_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper274_U0_fifo_w_out_V_V_write_pass_0_in = PE_wrapper274_U0_fifo_w_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_10_4_V_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_10_4_V_V_full_n_pass_1_q0 <= fifo_cin_PE_10_4_V_V_full_n_pass_1_out;
  end
  assign fifo_cin_PE_10_4_V_V_full_n_pass_1_in = fifo_cin_PE_10_4_V_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper226_U0_fifo_cin_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper226_U0_fifo_cin_out_V_V_din_pass_0_q0 <= PE_wrapper226_U0_fifo_cin_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper226_U0_fifo_cin_out_V_V_din_pass_0_in = PE_wrapper226_U0_fifo_cin_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper226_U0_fifo_cin_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper226_U0_fifo_cin_out_V_V_write_pass_0_q0 <= PE_wrapper226_U0_fifo_cin_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper226_U0_fifo_cin_out_V_V_write_pass_0_in = PE_wrapper226_U0_fifo_cin_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [31:0] PE_wrapper318_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper318_U0_fifo_cout_drain_out_V_din_pass_0_q0 <= PE_wrapper318_U0_fifo_cout_drain_out_V_din_pass_0_out;
  end
  assign PE_wrapper318_U0_fifo_cout_drain_out_V_din_pass_0_in = PE_wrapper318_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper318_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper318_U0_fifo_cout_drain_out_V_write_pass_0_q0 <= PE_wrapper318_U0_fifo_cout_drain_out_V_write_pass_0_out;
  end
  assign PE_wrapper318_U0_fifo_cout_drain_out_V_write_pass_0_in = PE_wrapper318_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [31:0] PE_wrapper274_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper274_U0_fifo_cout_drain_out_V_din_pass_0_q0 <= PE_wrapper274_U0_fifo_cout_drain_out_V_din_pass_0_out;
  end
  assign PE_wrapper274_U0_fifo_cout_drain_out_V_din_pass_0_in = PE_wrapper274_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper274_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper274_U0_fifo_cout_drain_out_V_write_pass_0_q0 <= PE_wrapper274_U0_fifo_cout_drain_out_V_write_pass_0_out;
  end
  assign PE_wrapper274_U0_fifo_cout_drain_out_V_write_pass_0_in = PE_wrapper274_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_PE_12_2_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_PE_12_2_V_full_n_pass_1_q0 <= fifo_cout_drain_PE_12_2_V_full_n_pass_1_out;
  end
  assign fifo_cout_drain_PE_12_2_V_full_n_pass_1_in = fifo_cout_drain_PE_12_2_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper321_U0_fifo_w_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper321_U0_fifo_w_out_V_V_din_pass_0_q0 <= PE_wrapper321_U0_fifo_w_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper321_U0_fifo_w_out_V_V_din_pass_0_in = PE_wrapper321_U0_fifo_w_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper321_U0_fifo_w_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper321_U0_fifo_w_out_V_V_write_pass_0_q0 <= PE_wrapper321_U0_fifo_w_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper321_U0_fifo_w_out_V_V_write_pass_0_in = PE_wrapper321_U0_fifo_w_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_PE_14_4_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_PE_14_4_V_full_n_pass_0_q0 <= fifo_cout_drain_PE_14_4_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_PE_14_4_V_full_n_pass_0_in = fifo_cout_drain_PE_14_4_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_cout_drain_IO_L1_out_2_13_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_cout_drain_IO_L1_out_2_13_V_V_full_n_pass_0_q0 <= fifo_cout_drain_cout_drain_IO_L1_out_2_13_V_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_cout_drain_IO_L1_out_2_13_V_V_full_n_pass_0_in = fifo_cout_drain_cout_drain_IO_L1_out_2_13_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg [63:0] cout_drain_IO_L1_out_wrapper434_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper434_U0_fifo_cout_drain_out_V_V_din_pass_0_q0 <= cout_drain_IO_L1_out_wrapper434_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper434_U0_fifo_cout_drain_out_V_V_din_pass_0_in = cout_drain_IO_L1_out_wrapper434_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  cout_drain_IO_L1_out_wrapper434_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper434_U0_fifo_cout_drain_out_V_V_write_pass_0_q0 <= cout_drain_IO_L1_out_wrapper434_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper434_U0_fifo_cout_drain_out_V_V_write_pass_0_in = cout_drain_IO_L1_out_wrapper434_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_PE_12_4_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_PE_12_4_V_full_n_pass_0_q0 <= fifo_cout_drain_PE_12_4_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_PE_12_4_V_full_n_pass_0_in = fifo_cout_drain_PE_12_4_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  ap_done_Boundary_X2Y6_To_X4Y6_q0;
  always @ (posedge ap_clk) begin
    ap_done_Boundary_X2Y6_To_X4Y6_q0 <= ap_done_Boundary_X2Y6_To_X4Y6_out;
  end
  assign ap_done_Boundary_X2Y6_To_X4Y6_in = ap_done_Boundary_X2Y6_To_X4Y6_q0;
  (* dont_touch = "yes" *) reg  ap_start_Boundary_X2Y8_To_X4Y8_q0;
  always @ (posedge ap_clk) begin
    ap_start_Boundary_X2Y8_To_X4Y8_q0 <= ap_start_Boundary_X2Y8_To_X4Y8_out;
  end
  assign ap_start_Boundary_X2Y8_To_X4Y8_in = ap_start_Boundary_X2Y8_To_X4Y8_q0;
  (* dont_touch = "yes" *) reg  ap_rst_n_Boundary_X2Y8_To_X4Y8_q0;
  always @ (posedge ap_clk) begin
    ap_rst_n_Boundary_X2Y8_To_X4Y8_q0 <= ap_rst_n_Boundary_X2Y8_To_X4Y8_out;
  end
  assign ap_rst_n_Boundary_X2Y8_To_X4Y8_in = ap_rst_n_Boundary_X2Y8_To_X4Y8_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper288_U0_fifo_cin_out_V_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper288_U0_fifo_cin_out_V_V_din_pass_1_q0 <= PE_wrapper288_U0_fifo_cin_out_V_V_din_pass_1_out;
  end
  assign PE_wrapper288_U0_fifo_cin_out_V_V_din_pass_1_in = PE_wrapper288_U0_fifo_cin_out_V_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_12_6_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_12_6_V_V_full_n_pass_0_q0 <= fifo_cin_PE_12_6_V_V_full_n_pass_0_out;
  end
  assign fifo_cin_PE_12_6_V_V_full_n_pass_0_in = fifo_cin_PE_12_6_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper288_U0_fifo_cin_out_V_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper288_U0_fifo_cin_out_V_V_write_pass_1_q0 <= PE_wrapper288_U0_fifo_cin_out_V_V_write_pass_1_out;
  end
  assign PE_wrapper288_U0_fifo_cin_out_V_V_write_pass_1_in = PE_wrapper288_U0_fifo_cin_out_V_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper311_U0_fifo_w_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper311_U0_fifo_w_out_V_V_din_pass_0_q0 <= PE_wrapper311_U0_fifo_w_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper311_U0_fifo_w_out_V_V_din_pass_0_in = PE_wrapper311_U0_fifo_w_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper311_U0_fifo_w_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper311_U0_fifo_w_out_V_V_write_pass_0_q0 <= PE_wrapper311_U0_fifo_w_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper311_U0_fifo_w_out_V_V_write_pass_0_in = PE_wrapper311_U0_fifo_w_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_9_5_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_9_5_V_V_full_n_pass_0_q0 <= fifo_cin_PE_9_5_V_V_full_n_pass_0_out;
  end
  assign fifo_cin_PE_9_5_V_V_full_n_pass_0_in = fifo_cin_PE_9_5_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper299_U0_fifo_w_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper299_U0_fifo_w_out_V_V_din_pass_0_q0 <= PE_wrapper299_U0_fifo_w_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper299_U0_fifo_w_out_V_V_din_pass_0_in = PE_wrapper299_U0_fifo_w_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper299_U0_fifo_w_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper299_U0_fifo_w_out_V_V_write_pass_0_q0 <= PE_wrapper299_U0_fifo_w_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper299_U0_fifo_w_out_V_V_write_pass_0_in = PE_wrapper299_U0_fifo_w_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [31:0] PE_wrapper263_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper263_U0_fifo_cout_drain_out_V_din_pass_0_q0 <= PE_wrapper263_U0_fifo_cout_drain_out_V_din_pass_0_out;
  end
  assign PE_wrapper263_U0_fifo_cout_drain_out_V_din_pass_0_in = PE_wrapper263_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper263_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper263_U0_fifo_cout_drain_out_V_write_pass_0_q0 <= PE_wrapper263_U0_fifo_cout_drain_out_V_write_pass_0_out;
  end
  assign PE_wrapper263_U0_fifo_cout_drain_out_V_write_pass_0_in = PE_wrapper263_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_13_5_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_13_5_V_V_full_n_pass_0_q0 <= fifo_w_PE_13_5_V_V_full_n_pass_0_out;
  end
  assign fifo_w_PE_13_5_V_V_full_n_pass_0_in = fifo_w_PE_13_5_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg [31:0] PE_wrapper336_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper336_U0_fifo_cout_drain_out_V_din_pass_0_q0 <= PE_wrapper336_U0_fifo_cout_drain_out_V_din_pass_0_out;
  end
  assign PE_wrapper336_U0_fifo_cout_drain_out_V_din_pass_0_in = PE_wrapper336_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper336_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper336_U0_fifo_cout_drain_out_V_write_pass_0_q0 <= PE_wrapper336_U0_fifo_cout_drain_out_V_write_pass_0_out;
  end
  assign PE_wrapper336_U0_fifo_cout_drain_out_V_write_pass_0_in = PE_wrapper336_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_9_5_V_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_9_5_V_V_full_n_pass_1_q0 <= fifo_w_PE_9_5_V_V_full_n_pass_1_out;
  end
  assign fifo_w_PE_9_5_V_V_full_n_pass_1_in = fifo_w_PE_9_5_V_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper337_U0_fifo_w_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper337_U0_fifo_w_out_V_V_din_pass_0_q0 <= PE_wrapper337_U0_fifo_w_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper337_U0_fifo_w_out_V_V_din_pass_0_in = PE_wrapper337_U0_fifo_w_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper337_U0_fifo_w_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper337_U0_fifo_w_out_V_V_write_pass_0_q0 <= PE_wrapper337_U0_fifo_w_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper337_U0_fifo_w_out_V_V_write_pass_0_in = PE_wrapper337_U0_fifo_w_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [63:0] cout_drain_IO_L1_out_wrapper450_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper450_U0_fifo_cout_drain_out_V_V_din_pass_0_q0 <= cout_drain_IO_L1_out_wrapper450_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper450_U0_fifo_cout_drain_out_V_V_din_pass_0_in = cout_drain_IO_L1_out_wrapper450_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  cout_drain_IO_L1_out_wrapper450_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper450_U0_fifo_cout_drain_out_V_V_write_pass_0_q0 <= cout_drain_IO_L1_out_wrapper450_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper450_U0_fifo_cout_drain_out_V_V_write_pass_0_in = cout_drain_IO_L1_out_wrapper450_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_12_5_V_V_full_n_pass_2_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_12_5_V_V_full_n_pass_2_q0 <= fifo_w_PE_12_5_V_V_full_n_pass_2_out;
  end
  assign fifo_w_PE_12_5_V_V_full_n_pass_2_in = fifo_w_PE_12_5_V_V_full_n_pass_2_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_14_5_V_V_full_n_pass_2_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_14_5_V_V_full_n_pass_2_q0 <= fifo_w_PE_14_5_V_V_full_n_pass_2_out;
  end
  assign fifo_w_PE_14_5_V_V_full_n_pass_2_in = fifo_w_PE_14_5_V_V_full_n_pass_2_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper263_U0_fifo_w_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper263_U0_fifo_w_out_V_V_din_pass_0_q0 <= PE_wrapper263_U0_fifo_w_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper263_U0_fifo_w_out_V_V_din_pass_0_in = PE_wrapper263_U0_fifo_w_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper263_U0_fifo_w_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper263_U0_fifo_w_out_V_V_write_pass_0_q0 <= PE_wrapper263_U0_fifo_w_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper263_U0_fifo_w_out_V_V_write_pass_0_in = PE_wrapper263_U0_fifo_w_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper323_U0_fifo_w_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper323_U0_fifo_w_out_V_V_din_pass_0_q0 <= PE_wrapper323_U0_fifo_w_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper323_U0_fifo_w_out_V_V_din_pass_0_in = PE_wrapper323_U0_fifo_w_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper323_U0_fifo_w_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper323_U0_fifo_w_out_V_V_write_pass_0_q0 <= PE_wrapper323_U0_fifo_w_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper323_U0_fifo_w_out_V_V_write_pass_0_in = PE_wrapper323_U0_fifo_w_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [31:0] PE_wrapper337_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper337_U0_fifo_cout_drain_out_V_din_pass_0_q0 <= PE_wrapper337_U0_fifo_cout_drain_out_V_din_pass_0_out;
  end
  assign PE_wrapper337_U0_fifo_cout_drain_out_V_din_pass_0_in = PE_wrapper337_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper337_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper337_U0_fifo_cout_drain_out_V_write_pass_0_q0 <= PE_wrapper337_U0_fifo_cout_drain_out_V_write_pass_0_out;
  end
  assign PE_wrapper337_U0_fifo_cout_drain_out_V_write_pass_0_in = PE_wrapper337_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_15_6_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_15_6_V_V_full_n_pass_0_q0 <= fifo_cin_PE_15_6_V_V_full_n_pass_0_out;
  end
  assign fifo_cin_PE_15_6_V_V_full_n_pass_0_in = fifo_cin_PE_15_6_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_15_5_V_V_full_n_pass_2_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_15_5_V_V_full_n_pass_2_q0 <= fifo_w_PE_15_5_V_V_full_n_pass_2_out;
  end
  assign fifo_w_PE_15_5_V_V_full_n_pass_2_in = fifo_w_PE_15_5_V_V_full_n_pass_2_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper263_U0_fifo_cin_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper263_U0_fifo_cin_out_V_V_din_pass_0_q0 <= PE_wrapper263_U0_fifo_cin_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper263_U0_fifo_cin_out_V_V_din_pass_0_in = PE_wrapper263_U0_fifo_cin_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper263_U0_fifo_cin_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper263_U0_fifo_cin_out_V_V_write_pass_0_q0 <= PE_wrapper263_U0_fifo_cin_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper263_U0_fifo_cin_out_V_V_write_pass_0_in = PE_wrapper263_U0_fifo_cin_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_15_7_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_15_7_V_V_full_n_pass_0_q0 <= fifo_cin_PE_15_7_V_V_full_n_pass_0_out;
  end
  assign fifo_cin_PE_15_7_V_V_full_n_pass_0_in = fifo_cin_PE_15_7_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_12_5_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_12_5_V_V_full_n_pass_0_q0 <= fifo_cin_PE_12_5_V_V_full_n_pass_0_out;
  end
  assign fifo_cin_PE_12_5_V_V_full_n_pass_0_in = fifo_cin_PE_12_5_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  ap_done_Boundary_X0Y8_To_X2Y8_q0;
  always @ (posedge ap_clk) begin
    ap_done_Boundary_X0Y8_To_X2Y8_q0 <= ap_done_Boundary_X0Y8_To_X2Y8_out;
  end
  assign ap_done_Boundary_X0Y8_To_X2Y8_in = ap_done_Boundary_X0Y8_To_X2Y8_q0;
  (* dont_touch = "yes" *) reg  ap_start_Boundary_X0Y10_To_X2Y10_q0;
  always @ (posedge ap_clk) begin
    ap_start_Boundary_X0Y10_To_X2Y10_q0 <= ap_start_Boundary_X0Y10_To_X2Y10_out;
  end
  assign ap_start_Boundary_X0Y10_To_X2Y10_in = ap_start_Boundary_X0Y10_To_X2Y10_q0;
  (* dont_touch = "yes" *) reg  ap_rst_n_Boundary_X0Y10_To_X2Y10_q0;
  always @ (posedge ap_clk) begin
    ap_rst_n_Boundary_X0Y10_To_X2Y10_q0 <= ap_rst_n_Boundary_X0Y10_To_X2Y10_out;
  end
  assign ap_rst_n_Boundary_X0Y10_To_X2Y10_in = ap_rst_n_Boundary_X0Y10_To_X2Y10_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper337_U0_fifo_w_out_V_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper337_U0_fifo_w_out_V_V_din_pass_1_q0 <= PE_wrapper337_U0_fifo_w_out_V_V_din_pass_1_out;
  end
  assign PE_wrapper337_U0_fifo_w_out_V_V_din_pass_1_in = PE_wrapper337_U0_fifo_w_out_V_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_15_8_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_15_8_V_V_full_n_pass_0_q0 <= fifo_w_PE_15_8_V_V_full_n_pass_0_out;
  end
  assign fifo_w_PE_15_8_V_V_full_n_pass_0_in = fifo_w_PE_15_8_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper337_U0_fifo_w_out_V_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper337_U0_fifo_w_out_V_V_write_pass_1_q0 <= PE_wrapper337_U0_fifo_w_out_V_V_write_pass_1_out;
  end
  assign PE_wrapper337_U0_fifo_w_out_V_V_write_pass_1_in = PE_wrapper337_U0_fifo_w_out_V_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_13_6_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_13_6_V_V_full_n_pass_0_q0 <= fifo_w_PE_13_6_V_V_full_n_pass_0_out;
  end
  assign fifo_w_PE_13_6_V_V_full_n_pass_0_in = fifo_w_PE_13_6_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_12_6_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_12_6_V_V_full_n_pass_0_q0 <= fifo_w_PE_12_6_V_V_full_n_pass_0_out;
  end
  assign fifo_w_PE_12_6_V_V_full_n_pass_0_in = fifo_w_PE_12_6_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_12_7_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_12_7_V_V_full_n_pass_0_q0 <= fifo_cin_PE_12_7_V_V_full_n_pass_0_out;
  end
  assign fifo_cin_PE_12_7_V_V_full_n_pass_0_in = fifo_cin_PE_12_7_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg [63:0] cout_drain_IO_L1_out_wrapper466_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper466_U0_fifo_cout_drain_out_V_V_din_pass_0_q0 <= cout_drain_IO_L1_out_wrapper466_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper466_U0_fifo_cout_drain_out_V_V_din_pass_0_in = cout_drain_IO_L1_out_wrapper466_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  cout_drain_IO_L1_out_wrapper466_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper466_U0_fifo_cout_drain_out_V_V_write_pass_0_q0 <= cout_drain_IO_L1_out_wrapper466_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper466_U0_fifo_cout_drain_out_V_V_write_pass_0_in = cout_drain_IO_L1_out_wrapper466_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_12_8_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_12_8_V_V_full_n_pass_0_q0 <= fifo_cin_PE_12_8_V_V_full_n_pass_0_out;
  end
  assign fifo_cin_PE_12_8_V_V_full_n_pass_0_in = fifo_cin_PE_12_8_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper302_U0_fifo_w_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper302_U0_fifo_w_out_V_V_din_pass_0_q0 <= PE_wrapper302_U0_fifo_w_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper302_U0_fifo_w_out_V_V_din_pass_0_in = PE_wrapper302_U0_fifo_w_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper302_U0_fifo_w_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper302_U0_fifo_w_out_V_V_write_pass_0_q0 <= PE_wrapper302_U0_fifo_w_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper302_U0_fifo_w_out_V_V_write_pass_0_in = PE_wrapper302_U0_fifo_w_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper325_U0_fifo_w_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper325_U0_fifo_w_out_V_V_din_pass_0_q0 <= PE_wrapper325_U0_fifo_w_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper325_U0_fifo_w_out_V_V_din_pass_0_in = PE_wrapper325_U0_fifo_w_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper325_U0_fifo_w_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper325_U0_fifo_w_out_V_V_write_pass_0_q0 <= PE_wrapper325_U0_fifo_w_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper325_U0_fifo_w_out_V_V_write_pass_0_in = PE_wrapper325_U0_fifo_w_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_PE_15_6_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_PE_15_6_V_full_n_pass_0_q0 <= fifo_cout_drain_PE_15_6_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_PE_15_6_V_full_n_pass_0_in = fifo_cout_drain_PE_15_6_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg [31:0] PE_wrapper302_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper302_U0_fifo_cout_drain_out_V_din_pass_0_q0 <= PE_wrapper302_U0_fifo_cout_drain_out_V_din_pass_0_out;
  end
  assign PE_wrapper302_U0_fifo_cout_drain_out_V_din_pass_0_in = PE_wrapper302_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper302_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper302_U0_fifo_cout_drain_out_V_write_pass_0_q0 <= PE_wrapper302_U0_fifo_cout_drain_out_V_write_pass_0_out;
  end
  assign PE_wrapper302_U0_fifo_cout_drain_out_V_write_pass_0_in = PE_wrapper302_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper302_U0_fifo_cin_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper302_U0_fifo_cin_out_V_V_din_pass_0_q0 <= PE_wrapper302_U0_fifo_cin_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper302_U0_fifo_cin_out_V_V_din_pass_0_in = PE_wrapper302_U0_fifo_cin_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper302_U0_fifo_cin_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper302_U0_fifo_cin_out_V_V_write_pass_0_q0 <= PE_wrapper302_U0_fifo_cin_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper302_U0_fifo_cin_out_V_V_write_pass_0_in = PE_wrapper302_U0_fifo_cin_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_12_6_V_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_12_6_V_V_full_n_pass_1_q0 <= fifo_cin_PE_12_6_V_V_full_n_pass_1_out;
  end
  assign fifo_cin_PE_12_6_V_V_full_n_pass_1_in = fifo_cin_PE_12_6_V_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_14_6_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_14_6_V_V_full_n_pass_0_q0 <= fifo_w_PE_14_6_V_V_full_n_pass_0_out;
  end
  assign fifo_w_PE_14_6_V_V_full_n_pass_0_in = fifo_w_PE_14_6_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_PE_15_7_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_PE_15_7_V_full_n_pass_0_q0 <= fifo_cout_drain_PE_15_7_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_PE_15_7_V_full_n_pass_0_in = fifo_cout_drain_PE_15_7_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper324_U0_fifo_cin_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper324_U0_fifo_cin_out_V_V_din_pass_0_q0 <= PE_wrapper324_U0_fifo_cin_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper324_U0_fifo_cin_out_V_V_din_pass_0_in = PE_wrapper324_U0_fifo_cin_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper324_U0_fifo_cin_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper324_U0_fifo_cin_out_V_V_write_pass_0_q0 <= PE_wrapper324_U0_fifo_cin_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper324_U0_fifo_cin_out_V_V_write_pass_0_in = PE_wrapper324_U0_fifo_cin_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper313_U0_fifo_w_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper313_U0_fifo_w_out_V_V_din_pass_0_q0 <= PE_wrapper313_U0_fifo_w_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper313_U0_fifo_w_out_V_V_din_pass_0_in = PE_wrapper313_U0_fifo_w_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper313_U0_fifo_w_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper313_U0_fifo_w_out_V_V_write_pass_0_q0 <= PE_wrapper313_U0_fifo_w_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper313_U0_fifo_w_out_V_V_write_pass_0_in = PE_wrapper313_U0_fifo_w_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper325_U0_fifo_cin_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper325_U0_fifo_cin_out_V_V_din_pass_0_q0 <= PE_wrapper325_U0_fifo_cin_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper325_U0_fifo_cin_out_V_V_din_pass_0_in = PE_wrapper325_U0_fifo_cin_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper325_U0_fifo_cin_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper325_U0_fifo_cin_out_V_V_write_pass_0_q0 <= PE_wrapper325_U0_fifo_cin_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper325_U0_fifo_cin_out_V_V_write_pass_0_in = PE_wrapper325_U0_fifo_cin_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [63:0] cout_drain_IO_L1_out_wrapper482_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper482_U0_fifo_cout_drain_out_V_V_din_pass_0_q0 <= cout_drain_IO_L1_out_wrapper482_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper482_U0_fifo_cout_drain_out_V_V_din_pass_0_in = cout_drain_IO_L1_out_wrapper482_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  cout_drain_IO_L1_out_wrapper482_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper482_U0_fifo_cout_drain_out_V_V_write_pass_0_q0 <= cout_drain_IO_L1_out_wrapper482_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper482_U0_fifo_cout_drain_out_V_V_write_pass_0_in = cout_drain_IO_L1_out_wrapper482_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  ap_done_Boundary_X0Y10_To_X2Y10_q0;
  always @ (posedge ap_clk) begin
    ap_done_Boundary_X0Y10_To_X2Y10_q0 <= ap_done_Boundary_X0Y10_To_X2Y10_out;
  end
  assign ap_done_Boundary_X0Y10_To_X2Y10_in = ap_done_Boundary_X0Y10_To_X2Y10_q0;
  (* dont_touch = "yes" *) reg  ap_start_Boundary_X0Y12_To_X2Y12_q0;
  always @ (posedge ap_clk) begin
    ap_start_Boundary_X0Y12_To_X2Y12_q0 <= ap_start_Boundary_X0Y12_To_X2Y12_out;
  end
  assign ap_start_Boundary_X0Y12_To_X2Y12_in = ap_start_Boundary_X0Y12_To_X2Y12_q0;
  (* dont_touch = "yes" *) reg  ap_rst_n_Boundary_X0Y12_To_X2Y12_q0;
  always @ (posedge ap_clk) begin
    ap_rst_n_Boundary_X0Y12_To_X2Y12_q0 <= ap_rst_n_Boundary_X0Y12_To_X2Y12_out;
  end
  assign ap_rst_n_Boundary_X0Y12_To_X2Y12_in = ap_rst_n_Boundary_X0Y12_To_X2Y12_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper263_U0_fifo_w_out_V_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper263_U0_fifo_w_out_V_V_din_pass_1_q0 <= PE_wrapper263_U0_fifo_w_out_V_V_din_pass_1_out;
  end
  assign PE_wrapper263_U0_fifo_w_out_V_V_din_pass_1_in = PE_wrapper263_U0_fifo_w_out_V_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_9_6_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_9_6_V_V_full_n_pass_0_q0 <= fifo_w_PE_9_6_V_V_full_n_pass_0_out;
  end
  assign fifo_w_PE_9_6_V_V_full_n_pass_0_in = fifo_w_PE_9_6_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper263_U0_fifo_w_out_V_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper263_U0_fifo_w_out_V_V_write_pass_1_q0 <= PE_wrapper263_U0_fifo_w_out_V_V_write_pass_1_out;
  end
  assign PE_wrapper263_U0_fifo_w_out_V_V_write_pass_1_in = PE_wrapper263_U0_fifo_w_out_V_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper251_U0_fifo_cin_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper251_U0_fifo_cin_out_V_V_din_pass_0_q0 <= PE_wrapper251_U0_fifo_cin_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper251_U0_fifo_cin_out_V_V_din_pass_0_in = PE_wrapper251_U0_fifo_cin_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper251_U0_fifo_cin_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper251_U0_fifo_cin_out_V_V_write_pass_0_q0 <= PE_wrapper251_U0_fifo_cin_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper251_U0_fifo_cin_out_V_V_write_pass_0_in = PE_wrapper251_U0_fifo_cin_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_PE_9_5_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_PE_9_5_V_full_n_pass_0_q0 <= fifo_cout_drain_PE_9_5_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_PE_9_5_V_full_n_pass_0_in = fifo_cout_drain_PE_9_5_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper276_U0_fifo_w_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper276_U0_fifo_w_out_V_V_din_pass_0_q0 <= PE_wrapper276_U0_fifo_w_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper276_U0_fifo_w_out_V_V_din_pass_0_in = PE_wrapper276_U0_fifo_w_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper276_U0_fifo_w_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper276_U0_fifo_w_out_V_V_write_pass_0_q0 <= PE_wrapper276_U0_fifo_w_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper276_U0_fifo_w_out_V_V_write_pass_0_in = PE_wrapper276_U0_fifo_w_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_PE_9_6_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_PE_9_6_V_full_n_pass_0_q0 <= fifo_cout_drain_PE_9_6_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_PE_9_6_V_full_n_pass_0_in = fifo_cout_drain_PE_9_6_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_cout_drain_IO_L1_out_6_12_V_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_cout_drain_IO_L1_out_6_12_V_V_full_n_pass_1_q0 <= fifo_cout_drain_cout_drain_IO_L1_out_6_12_V_V_full_n_pass_1_out;
  end
  assign fifo_cout_drain_cout_drain_IO_L1_out_6_12_V_V_full_n_pass_1_in = fifo_cout_drain_cout_drain_IO_L1_out_6_12_V_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_10_6_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_10_6_V_V_full_n_pass_0_q0 <= fifo_cin_PE_10_6_V_V_full_n_pass_0_out;
  end
  assign fifo_cin_PE_10_6_V_V_full_n_pass_0_in = fifo_cin_PE_10_6_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_11_5_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_11_5_V_V_full_n_pass_0_q0 <= fifo_w_PE_11_5_V_V_full_n_pass_0_out;
  end
  assign fifo_w_PE_11_5_V_V_full_n_pass_0_in = fifo_w_PE_11_5_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_6_5_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_6_5_V_V_full_n_pass_0_q0 <= fifo_cin_PE_6_5_V_V_full_n_pass_0_out;
  end
  assign fifo_cin_PE_6_5_V_V_full_n_pass_0_in = fifo_cin_PE_6_5_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper227_U0_fifo_w_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper227_U0_fifo_w_out_V_V_din_pass_0_q0 <= PE_wrapper227_U0_fifo_w_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper227_U0_fifo_w_out_V_V_din_pass_0_in = PE_wrapper227_U0_fifo_w_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper227_U0_fifo_w_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper227_U0_fifo_w_out_V_V_write_pass_0_q0 <= PE_wrapper227_U0_fifo_w_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper227_U0_fifo_w_out_V_V_write_pass_0_in = PE_wrapper227_U0_fifo_w_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_8_5_V_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_8_5_V_V_full_n_pass_1_q0 <= fifo_w_PE_8_5_V_V_full_n_pass_1_out;
  end
  assign fifo_w_PE_8_5_V_V_full_n_pass_1_in = fifo_w_PE_8_5_V_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_cout_drain_IO_L1_out_5_12_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_cout_drain_IO_L1_out_5_12_V_V_full_n_pass_0_q0 <= fifo_cout_drain_cout_drain_IO_L1_out_5_12_V_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_cout_drain_IO_L1_out_5_12_V_V_full_n_pass_0_in = fifo_cout_drain_cout_drain_IO_L1_out_5_12_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_6_5_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_6_5_V_V_full_n_pass_0_q0 <= fifo_w_PE_6_5_V_V_full_n_pass_0_out;
  end
  assign fifo_w_PE_6_5_V_V_full_n_pass_0_in = fifo_w_PE_6_5_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg [63:0] cout_drain_IO_L1_out_wrapper456_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper456_U0_fifo_cout_drain_out_V_V_din_pass_0_q0 <= cout_drain_IO_L1_out_wrapper456_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper456_U0_fifo_cout_drain_out_V_V_din_pass_0_in = cout_drain_IO_L1_out_wrapper456_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  cout_drain_IO_L1_out_wrapper456_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper456_U0_fifo_cout_drain_out_V_V_write_pass_0_q0 <= cout_drain_IO_L1_out_wrapper456_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper456_U0_fifo_cout_drain_out_V_V_write_pass_0_in = cout_drain_IO_L1_out_wrapper456_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper288_U0_fifo_cin_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper288_U0_fifo_cin_out_V_V_din_pass_0_q0 <= PE_wrapper288_U0_fifo_cin_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper288_U0_fifo_cin_out_V_V_din_pass_0_in = PE_wrapper288_U0_fifo_cin_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper288_U0_fifo_cin_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper288_U0_fifo_cin_out_V_V_write_pass_0_q0 <= PE_wrapper288_U0_fifo_cin_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper288_U0_fifo_cin_out_V_V_write_pass_0_in = PE_wrapper288_U0_fifo_cin_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper251_U0_fifo_w_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper251_U0_fifo_w_out_V_V_din_pass_0_q0 <= PE_wrapper251_U0_fifo_w_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper251_U0_fifo_w_out_V_V_din_pass_0_in = PE_wrapper251_U0_fifo_w_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper251_U0_fifo_w_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper251_U0_fifo_w_out_V_V_write_pass_0_q0 <= PE_wrapper251_U0_fifo_w_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper251_U0_fifo_w_out_V_V_write_pass_0_in = PE_wrapper251_U0_fifo_w_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_10_5_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_10_5_V_V_full_n_pass_0_q0 <= fifo_w_PE_10_5_V_V_full_n_pass_0_out;
  end
  assign fifo_w_PE_10_5_V_V_full_n_pass_0_in = fifo_w_PE_10_5_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper239_U0_fifo_w_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper239_U0_fifo_w_out_V_V_din_pass_0_q0 <= PE_wrapper239_U0_fifo_w_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper239_U0_fifo_w_out_V_V_din_pass_0_in = PE_wrapper239_U0_fifo_w_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper239_U0_fifo_w_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper239_U0_fifo_w_out_V_V_write_pass_0_q0 <= PE_wrapper239_U0_fifo_w_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper239_U0_fifo_w_out_V_V_write_pass_0_in = PE_wrapper239_U0_fifo_w_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_7_5_V_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_7_5_V_V_full_n_pass_1_q0 <= fifo_w_PE_7_5_V_V_full_n_pass_1_out;
  end
  assign fifo_w_PE_7_5_V_V_full_n_pass_1_in = fifo_w_PE_7_5_V_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_10_5_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_10_5_V_V_full_n_pass_0_q0 <= fifo_cin_PE_10_5_V_V_full_n_pass_0_out;
  end
  assign fifo_cin_PE_10_5_V_V_full_n_pass_0_in = fifo_cin_PE_10_5_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg [63:0] cout_drain_IO_L1_out_wrapper469_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper469_U0_fifo_cout_drain_out_V_V_din_pass_0_q0 <= cout_drain_IO_L1_out_wrapper469_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper469_U0_fifo_cout_drain_out_V_V_din_pass_0_in = cout_drain_IO_L1_out_wrapper469_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  cout_drain_IO_L1_out_wrapper469_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper469_U0_fifo_cout_drain_out_V_V_write_pass_0_q0 <= cout_drain_IO_L1_out_wrapper469_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper469_U0_fifo_cout_drain_out_V_V_write_pass_0_in = cout_drain_IO_L1_out_wrapper469_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper288_U0_fifo_w_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper288_U0_fifo_w_out_V_V_din_pass_0_q0 <= PE_wrapper288_U0_fifo_w_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper288_U0_fifo_w_out_V_V_din_pass_0_in = PE_wrapper288_U0_fifo_w_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper288_U0_fifo_w_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper288_U0_fifo_w_out_V_V_write_pass_0_q0 <= PE_wrapper288_U0_fifo_w_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper288_U0_fifo_w_out_V_V_write_pass_0_in = PE_wrapper288_U0_fifo_w_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper287_U0_fifo_cin_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper287_U0_fifo_cin_out_V_V_din_pass_0_q0 <= PE_wrapper287_U0_fifo_cin_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper287_U0_fifo_cin_out_V_V_din_pass_0_in = PE_wrapper287_U0_fifo_cin_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper287_U0_fifo_cin_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper287_U0_fifo_cin_out_V_V_write_pass_0_q0 <= PE_wrapper287_U0_fifo_cin_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper287_U0_fifo_cin_out_V_V_write_pass_0_in = PE_wrapper287_U0_fifo_cin_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  ap_done_Boundary_X2Y8_To_X4Y8_q0;
  always @ (posedge ap_clk) begin
    ap_done_Boundary_X2Y8_To_X4Y8_q0 <= ap_done_Boundary_X2Y8_To_X4Y8_out;
  end
  assign ap_done_Boundary_X2Y8_To_X4Y8_in = ap_done_Boundary_X2Y8_To_X4Y8_q0;
  (* dont_touch = "yes" *) reg  ap_start_Boundary_X2Y10_To_X4Y10_q0;
  always @ (posedge ap_clk) begin
    ap_start_Boundary_X2Y10_To_X4Y10_q0 <= ap_start_Boundary_X2Y10_To_X4Y10_out;
  end
  assign ap_start_Boundary_X2Y10_To_X4Y10_in = ap_start_Boundary_X2Y10_To_X4Y10_q0;
  (* dont_touch = "yes" *) reg  ap_rst_n_Boundary_X2Y10_To_X4Y10_q0;
  always @ (posedge ap_clk) begin
    ap_rst_n_Boundary_X2Y10_To_X4Y10_q0 <= ap_rst_n_Boundary_X2Y10_To_X4Y10_out;
  end
  assign ap_rst_n_Boundary_X2Y10_To_X4Y10_in = ap_rst_n_Boundary_X2Y10_To_X4Y10_q0;
  (* dont_touch = "yes" *) reg [63:0] cout_drain_IO_L1_out_wrapper466_U0_fifo_cout_drain_out_V_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper466_U0_fifo_cout_drain_out_V_V_din_pass_1_q0 <= cout_drain_IO_L1_out_wrapper466_U0_fifo_cout_drain_out_V_V_din_pass_1_out;
  end
  assign cout_drain_IO_L1_out_wrapper466_U0_fifo_cout_drain_out_V_V_din_pass_1_in = cout_drain_IO_L1_out_wrapper466_U0_fifo_cout_drain_out_V_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_cout_drain_IO_L1_out_6_12_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_cout_drain_IO_L1_out_6_12_V_V_full_n_pass_0_q0 <= fifo_cout_drain_cout_drain_IO_L1_out_6_12_V_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_cout_drain_IO_L1_out_6_12_V_V_full_n_pass_0_in = fifo_cout_drain_cout_drain_IO_L1_out_6_12_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  cout_drain_IO_L1_out_wrapper466_U0_fifo_cout_drain_out_V_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper466_U0_fifo_cout_drain_out_V_V_write_pass_1_q0 <= cout_drain_IO_L1_out_wrapper466_U0_fifo_cout_drain_out_V_V_write_pass_1_out;
  end
  assign cout_drain_IO_L1_out_wrapper466_U0_fifo_cout_drain_out_V_V_write_pass_1_in = cout_drain_IO_L1_out_wrapper466_U0_fifo_cout_drain_out_V_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper302_U0_fifo_w_out_V_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper302_U0_fifo_w_out_V_V_din_pass_1_q0 <= PE_wrapper302_U0_fifo_w_out_V_V_din_pass_1_out;
  end
  assign PE_wrapper302_U0_fifo_w_out_V_V_din_pass_1_in = PE_wrapper302_U0_fifo_w_out_V_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_12_9_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_12_9_V_V_full_n_pass_0_q0 <= fifo_w_PE_12_9_V_V_full_n_pass_0_out;
  end
  assign fifo_w_PE_12_9_V_V_full_n_pass_0_in = fifo_w_PE_12_9_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper302_U0_fifo_w_out_V_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper302_U0_fifo_w_out_V_V_write_pass_1_q0 <= PE_wrapper302_U0_fifo_w_out_V_V_write_pass_1_out;
  end
  assign PE_wrapper302_U0_fifo_w_out_V_V_write_pass_1_in = PE_wrapper302_U0_fifo_w_out_V_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper290_U0_fifo_w_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper290_U0_fifo_w_out_V_V_din_pass_0_q0 <= PE_wrapper290_U0_fifo_w_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper290_U0_fifo_w_out_V_V_din_pass_0_in = PE_wrapper290_U0_fifo_w_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper290_U0_fifo_w_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper290_U0_fifo_w_out_V_V_write_pass_0_q0 <= PE_wrapper290_U0_fifo_w_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper290_U0_fifo_w_out_V_V_write_pass_0_in = PE_wrapper290_U0_fifo_w_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_9_7_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_9_7_V_V_full_n_pass_0_q0 <= fifo_cin_PE_9_7_V_V_full_n_pass_0_out;
  end
  assign fifo_cin_PE_9_7_V_V_full_n_pass_0_in = fifo_cin_PE_9_7_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper289_U0_fifo_cin_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper289_U0_fifo_cin_out_V_V_din_pass_0_q0 <= PE_wrapper289_U0_fifo_cin_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper289_U0_fifo_cin_out_V_V_din_pass_0_in = PE_wrapper289_U0_fifo_cin_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper289_U0_fifo_cin_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper289_U0_fifo_cin_out_V_V_write_pass_0_q0 <= PE_wrapper289_U0_fifo_cin_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper289_U0_fifo_cin_out_V_V_write_pass_0_in = PE_wrapper289_U0_fifo_cin_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_cout_drain_IO_L1_out_7_12_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_cout_drain_IO_L1_out_7_12_V_V_full_n_pass_0_q0 <= fifo_cout_drain_cout_drain_IO_L1_out_7_12_V_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_cout_drain_IO_L1_out_7_12_V_V_full_n_pass_0_in = fifo_cout_drain_cout_drain_IO_L1_out_7_12_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_10_7_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_10_7_V_V_full_n_pass_0_q0 <= fifo_w_PE_10_7_V_V_full_n_pass_0_out;
  end
  assign fifo_w_PE_10_7_V_V_full_n_pass_0_in = fifo_w_PE_10_7_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg [31:0] PE_wrapper264_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper264_U0_fifo_cout_drain_out_V_din_pass_0_q0 <= PE_wrapper264_U0_fifo_cout_drain_out_V_din_pass_0_out;
  end
  assign PE_wrapper264_U0_fifo_cout_drain_out_V_din_pass_0_in = PE_wrapper264_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper264_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper264_U0_fifo_cout_drain_out_V_write_pass_0_q0 <= PE_wrapper264_U0_fifo_cout_drain_out_V_write_pass_0_out;
  end
  assign PE_wrapper264_U0_fifo_cout_drain_out_V_write_pass_0_in = PE_wrapper264_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper278_U0_fifo_w_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper278_U0_fifo_w_out_V_V_din_pass_0_q0 <= PE_wrapper278_U0_fifo_w_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper278_U0_fifo_w_out_V_V_din_pass_0_in = PE_wrapper278_U0_fifo_w_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper278_U0_fifo_w_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper278_U0_fifo_w_out_V_V_write_pass_0_q0 <= PE_wrapper278_U0_fifo_w_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper278_U0_fifo_w_out_V_V_write_pass_0_in = PE_wrapper278_U0_fifo_w_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper290_U0_fifo_cin_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper290_U0_fifo_cin_out_V_V_din_pass_0_q0 <= PE_wrapper290_U0_fifo_cin_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper290_U0_fifo_cin_out_V_V_din_pass_0_in = PE_wrapper290_U0_fifo_cin_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper290_U0_fifo_cin_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper290_U0_fifo_cin_out_V_V_write_pass_0_q0 <= PE_wrapper290_U0_fifo_cin_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper290_U0_fifo_cin_out_V_V_write_pass_0_in = PE_wrapper290_U0_fifo_cin_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_cout_drain_IO_L1_out_8_13_V_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_cout_drain_IO_L1_out_8_13_V_V_full_n_pass_1_q0 <= fifo_cout_drain_cout_drain_IO_L1_out_8_13_V_V_full_n_pass_1_out;
  end
  assign fifo_cout_drain_cout_drain_IO_L1_out_8_13_V_V_full_n_pass_1_in = fifo_cout_drain_cout_drain_IO_L1_out_8_13_V_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper264_U0_fifo_cin_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper264_U0_fifo_cin_out_V_V_din_pass_0_q0 <= PE_wrapper264_U0_fifo_cin_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper264_U0_fifo_cin_out_V_V_din_pass_0_in = PE_wrapper264_U0_fifo_cin_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper264_U0_fifo_cin_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper264_U0_fifo_cin_out_V_V_write_pass_0_q0 <= PE_wrapper264_U0_fifo_cin_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper264_U0_fifo_cin_out_V_V_write_pass_0_in = PE_wrapper264_U0_fifo_cin_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_9_6_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_9_6_V_V_full_n_pass_0_q0 <= fifo_cin_PE_9_6_V_V_full_n_pass_0_out;
  end
  assign fifo_cin_PE_9_6_V_V_full_n_pass_0_in = fifo_cin_PE_9_6_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_PE_12_8_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_PE_12_8_V_full_n_pass_0_q0 <= fifo_cout_drain_PE_12_8_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_PE_12_8_V_full_n_pass_0_in = fifo_cout_drain_PE_12_8_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper266_U0_fifo_w_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper266_U0_fifo_w_out_V_V_din_pass_0_q0 <= PE_wrapper266_U0_fifo_w_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper266_U0_fifo_w_out_V_V_din_pass_0_in = PE_wrapper266_U0_fifo_w_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper266_U0_fifo_w_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper266_U0_fifo_w_out_V_V_write_pass_0_q0 <= PE_wrapper266_U0_fifo_w_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper266_U0_fifo_w_out_V_V_write_pass_0_in = PE_wrapper266_U0_fifo_w_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [63:0] cout_drain_IO_L1_out_wrapper501_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper501_U0_fifo_cout_drain_out_V_V_din_pass_0_q0 <= cout_drain_IO_L1_out_wrapper501_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper501_U0_fifo_cout_drain_out_V_V_din_pass_0_in = cout_drain_IO_L1_out_wrapper501_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  cout_drain_IO_L1_out_wrapper501_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper501_U0_fifo_cout_drain_out_V_V_write_pass_0_q0 <= cout_drain_IO_L1_out_wrapper501_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper501_U0_fifo_cout_drain_out_V_V_write_pass_0_in = cout_drain_IO_L1_out_wrapper501_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_9_6_V_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_9_6_V_V_full_n_pass_1_q0 <= fifo_w_PE_9_6_V_V_full_n_pass_1_out;
  end
  assign fifo_w_PE_9_6_V_V_full_n_pass_1_in = fifo_w_PE_9_6_V_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg [63:0] cout_drain_IO_L1_out_wrapper485_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper485_U0_fifo_cout_drain_out_V_V_din_pass_0_q0 <= cout_drain_IO_L1_out_wrapper485_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper485_U0_fifo_cout_drain_out_V_V_din_pass_0_in = cout_drain_IO_L1_out_wrapper485_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  cout_drain_IO_L1_out_wrapper485_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper485_U0_fifo_cout_drain_out_V_V_write_pass_0_q0 <= cout_drain_IO_L1_out_wrapper485_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper485_U0_fifo_cout_drain_out_V_V_write_pass_0_in = cout_drain_IO_L1_out_wrapper485_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_9_8_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_9_8_V_V_full_n_pass_0_q0 <= fifo_cin_PE_9_8_V_V_full_n_pass_0_out;
  end
  assign fifo_cin_PE_9_8_V_V_full_n_pass_0_in = fifo_cin_PE_9_8_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_11_7_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_11_7_V_V_full_n_pass_0_q0 <= fifo_w_PE_11_7_V_V_full_n_pass_0_out;
  end
  assign fifo_w_PE_11_7_V_V_full_n_pass_0_in = fifo_w_PE_11_7_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  ap_done_Boundary_X2Y10_To_X4Y10_q0;
  always @ (posedge ap_clk) begin
    ap_done_Boundary_X2Y10_To_X4Y10_q0 <= ap_done_Boundary_X2Y10_To_X4Y10_out;
  end
  assign ap_done_Boundary_X2Y10_To_X4Y10_in = ap_done_Boundary_X2Y10_To_X4Y10_q0;
  (* dont_touch = "yes" *) reg  ap_start_Boundary_X2Y12_To_X4Y12_q0;
  always @ (posedge ap_clk) begin
    ap_start_Boundary_X2Y12_To_X4Y12_q0 <= ap_start_Boundary_X2Y12_To_X4Y12_out;
  end
  assign ap_start_Boundary_X2Y12_To_X4Y12_in = ap_start_Boundary_X2Y12_To_X4Y12_q0;
  (* dont_touch = "yes" *) reg  ap_rst_n_Boundary_X2Y12_To_X4Y12_q0;
  always @ (posedge ap_clk) begin
    ap_rst_n_Boundary_X2Y12_To_X4Y12_q0 <= ap_rst_n_Boundary_X2Y12_To_X4Y12_out;
  end
  assign ap_rst_n_Boundary_X2Y12_To_X4Y12_in = ap_rst_n_Boundary_X2Y12_To_X4Y12_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper304_U0_fifo_cin_out_V_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper304_U0_fifo_cin_out_V_V_din_pass_1_q0 <= PE_wrapper304_U0_fifo_cin_out_V_V_din_pass_1_out;
  end
  assign PE_wrapper304_U0_fifo_cin_out_V_V_din_pass_1_in = PE_wrapper304_U0_fifo_cin_out_V_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_13_10_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_13_10_V_V_full_n_pass_0_q0 <= fifo_cin_PE_13_10_V_V_full_n_pass_0_out;
  end
  assign fifo_cin_PE_13_10_V_V_full_n_pass_0_in = fifo_cin_PE_13_10_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper304_U0_fifo_cin_out_V_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper304_U0_fifo_cin_out_V_V_write_pass_1_q0 <= PE_wrapper304_U0_fifo_cin_out_V_V_write_pass_1_out;
  end
  assign PE_wrapper304_U0_fifo_cin_out_V_V_write_pass_1_in = PE_wrapper304_U0_fifo_cin_out_V_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper305_U0_fifo_cin_out_V_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper305_U0_fifo_cin_out_V_V_din_pass_1_q0 <= PE_wrapper305_U0_fifo_cin_out_V_V_din_pass_1_out;
  end
  assign PE_wrapper305_U0_fifo_cin_out_V_V_din_pass_1_in = PE_wrapper305_U0_fifo_cin_out_V_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_13_11_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_13_11_V_V_full_n_pass_0_q0 <= fifo_cin_PE_13_11_V_V_full_n_pass_0_out;
  end
  assign fifo_cin_PE_13_11_V_V_full_n_pass_0_in = fifo_cin_PE_13_11_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper305_U0_fifo_cin_out_V_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper305_U0_fifo_cin_out_V_V_write_pass_1_q0 <= PE_wrapper305_U0_fifo_cin_out_V_V_write_pass_1_out;
  end
  assign PE_wrapper305_U0_fifo_cin_out_V_V_write_pass_1_in = PE_wrapper305_U0_fifo_cin_out_V_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [63:0] cout_drain_IO_L1_out_wrapper513_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper513_U0_fifo_cout_drain_out_V_V_din_pass_0_q0 <= cout_drain_IO_L1_out_wrapper513_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper513_U0_fifo_cout_drain_out_V_V_din_pass_0_in = cout_drain_IO_L1_out_wrapper513_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  cout_drain_IO_L1_out_wrapper513_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper513_U0_fifo_cout_drain_out_V_V_write_pass_0_q0 <= cout_drain_IO_L1_out_wrapper513_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper513_U0_fifo_cout_drain_out_V_V_write_pass_0_in = cout_drain_IO_L1_out_wrapper513_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_13_9_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_13_9_V_V_full_n_pass_0_q0 <= fifo_cin_PE_13_9_V_V_full_n_pass_0_out;
  end
  assign fifo_cin_PE_13_9_V_V_full_n_pass_0_in = fifo_cin_PE_13_9_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper327_U0_fifo_w_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper327_U0_fifo_w_out_V_V_din_pass_0_q0 <= PE_wrapper327_U0_fifo_w_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper327_U0_fifo_w_out_V_V_din_pass_0_in = PE_wrapper327_U0_fifo_w_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper327_U0_fifo_w_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper327_U0_fifo_w_out_V_V_write_pass_0_q0 <= PE_wrapper327_U0_fifo_w_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper327_U0_fifo_w_out_V_V_write_pass_0_in = PE_wrapper327_U0_fifo_w_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [63:0] cout_drain_IO_L1_out_wrapper497_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper497_U0_fifo_cout_drain_out_V_V_din_pass_0_q0 <= cout_drain_IO_L1_out_wrapper497_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper497_U0_fifo_cout_drain_out_V_V_din_pass_0_in = cout_drain_IO_L1_out_wrapper497_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  cout_drain_IO_L1_out_wrapper497_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper497_U0_fifo_cout_drain_out_V_V_write_pass_0_q0 <= cout_drain_IO_L1_out_wrapper497_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper497_U0_fifo_cout_drain_out_V_V_write_pass_0_in = cout_drain_IO_L1_out_wrapper497_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_14_8_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_14_8_V_V_full_n_pass_0_q0 <= fifo_w_PE_14_8_V_V_full_n_pass_0_out;
  end
  assign fifo_w_PE_14_8_V_V_full_n_pass_0_in = fifo_w_PE_14_8_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper315_U0_fifo_w_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper315_U0_fifo_w_out_V_V_din_pass_0_q0 <= PE_wrapper315_U0_fifo_w_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper315_U0_fifo_w_out_V_V_din_pass_0_in = PE_wrapper315_U0_fifo_w_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper315_U0_fifo_w_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper315_U0_fifo_w_out_V_V_write_pass_0_q0 <= PE_wrapper315_U0_fifo_w_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper315_U0_fifo_w_out_V_V_write_pass_0_in = PE_wrapper315_U0_fifo_w_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_13_8_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_13_8_V_V_full_n_pass_0_q0 <= fifo_cin_PE_13_8_V_V_full_n_pass_0_out;
  end
  assign fifo_cin_PE_13_8_V_V_full_n_pass_0_in = fifo_cin_PE_13_8_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_15_8_V_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_15_8_V_V_full_n_pass_1_q0 <= fifo_w_PE_15_8_V_V_full_n_pass_1_out;
  end
  assign fifo_w_PE_15_8_V_V_full_n_pass_1_in = fifo_w_PE_15_8_V_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_13_8_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_13_8_V_V_full_n_pass_0_q0 <= fifo_w_PE_13_8_V_V_full_n_pass_0_out;
  end
  assign fifo_w_PE_13_8_V_V_full_n_pass_0_in = fifo_w_PE_13_8_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper339_U0_fifo_w_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper339_U0_fifo_w_out_V_V_din_pass_0_q0 <= PE_wrapper339_U0_fifo_w_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper339_U0_fifo_w_out_V_V_din_pass_0_in = PE_wrapper339_U0_fifo_w_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper339_U0_fifo_w_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper339_U0_fifo_w_out_V_V_write_pass_0_q0 <= PE_wrapper339_U0_fifo_w_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper339_U0_fifo_w_out_V_V_write_pass_0_in = PE_wrapper339_U0_fifo_w_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  ap_done_Boundary_X0Y12_To_X2Y12_q0;
  always @ (posedge ap_clk) begin
    ap_done_Boundary_X0Y12_To_X2Y12_q0 <= ap_done_Boundary_X0Y12_To_X2Y12_out;
  end
  assign ap_done_Boundary_X0Y12_To_X2Y12_in = ap_done_Boundary_X0Y12_To_X2Y12_q0;
  (* dont_touch = "yes" *) reg  ap_start_Boundary_X0Y14_To_X2Y14_q0;
  always @ (posedge ap_clk) begin
    ap_start_Boundary_X0Y14_To_X2Y14_q0 <= ap_start_Boundary_X0Y14_To_X2Y14_out;
  end
  assign ap_start_Boundary_X0Y14_To_X2Y14_in = ap_start_Boundary_X0Y14_To_X2Y14_q0;
  (* dont_touch = "yes" *) reg  ap_rst_n_Boundary_X0Y14_To_X2Y14_q0;
  always @ (posedge ap_clk) begin
    ap_rst_n_Boundary_X0Y14_To_X2Y14_q0 <= ap_rst_n_Boundary_X0Y14_To_X2Y14_out;
  end
  assign ap_rst_n_Boundary_X0Y14_To_X2Y14_in = ap_rst_n_Boundary_X0Y14_To_X2Y14_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_13_10_V_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_13_10_V_V_full_n_pass_1_q0 <= fifo_cin_PE_13_10_V_V_full_n_pass_1_out;
  end
  assign fifo_cin_PE_13_10_V_V_full_n_pass_1_in = fifo_cin_PE_13_10_V_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_14_10_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_14_10_V_V_full_n_pass_0_q0 <= fifo_w_PE_14_10_V_V_full_n_pass_0_out;
  end
  assign fifo_w_PE_14_10_V_V_full_n_pass_0_in = fifo_w_PE_14_10_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_13_10_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_13_10_V_V_full_n_pass_0_q0 <= fifo_w_PE_13_10_V_V_full_n_pass_0_out;
  end
  assign fifo_w_PE_13_10_V_V_full_n_pass_0_in = fifo_w_PE_13_10_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg [63:0] cout_drain_IO_L1_out_wrapper529_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper529_U0_fifo_cout_drain_out_V_V_din_pass_0_q0 <= cout_drain_IO_L1_out_wrapper529_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper529_U0_fifo_cout_drain_out_V_V_din_pass_0_in = cout_drain_IO_L1_out_wrapper529_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  cout_drain_IO_L1_out_wrapper529_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper529_U0_fifo_cout_drain_out_V_V_write_pass_0_q0 <= cout_drain_IO_L1_out_wrapper529_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper529_U0_fifo_cout_drain_out_V_V_write_pass_0_in = cout_drain_IO_L1_out_wrapper529_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_13_11_V_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_13_11_V_V_full_n_pass_1_q0 <= fifo_cin_PE_13_11_V_V_full_n_pass_1_out;
  end
  assign fifo_cin_PE_13_11_V_V_full_n_pass_1_in = fifo_cin_PE_13_11_V_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_15_10_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_15_10_V_V_full_n_pass_0_q0 <= fifo_w_PE_15_10_V_V_full_n_pass_0_out;
  end
  assign fifo_w_PE_15_10_V_V_full_n_pass_0_in = fifo_w_PE_15_10_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg [63:0] cout_drain_IO_L1_out_wrapper544_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper544_U0_fifo_cout_drain_out_V_V_din_pass_0_q0 <= cout_drain_IO_L1_out_wrapper544_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper544_U0_fifo_cout_drain_out_V_V_din_pass_0_in = cout_drain_IO_L1_out_wrapper544_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  cout_drain_IO_L1_out_wrapper544_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper544_U0_fifo_cout_drain_out_V_V_write_pass_0_q0 <= cout_drain_IO_L1_out_wrapper544_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper544_U0_fifo_cout_drain_out_V_V_write_pass_0_in = cout_drain_IO_L1_out_wrapper544_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  ap_done_Boundary_X0Y14_To_X2Y14_q0;
  always @ (posedge ap_clk) begin
    ap_done_Boundary_X0Y14_To_X2Y14_q0 <= ap_done_Boundary_X0Y14_To_X2Y14_out;
  end
  assign ap_done_Boundary_X0Y14_To_X2Y14_in = ap_done_Boundary_X0Y14_To_X2Y14_q0;
  (* dont_touch = "yes" *) reg [63:0] cout_drain_IO_L1_out_wrapper497_U0_fifo_cout_drain_out_V_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper497_U0_fifo_cout_drain_out_V_V_din_pass_1_q0 <= cout_drain_IO_L1_out_wrapper497_U0_fifo_cout_drain_out_V_V_din_pass_1_out;
  end
  assign cout_drain_IO_L1_out_wrapper497_U0_fifo_cout_drain_out_V_V_din_pass_1_in = cout_drain_IO_L1_out_wrapper497_U0_fifo_cout_drain_out_V_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_cout_drain_IO_L1_out_8_13_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_cout_drain_IO_L1_out_8_13_V_V_full_n_pass_0_q0 <= fifo_cout_drain_cout_drain_IO_L1_out_8_13_V_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_cout_drain_IO_L1_out_8_13_V_V_full_n_pass_0_in = fifo_cout_drain_cout_drain_IO_L1_out_8_13_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  cout_drain_IO_L1_out_wrapper497_U0_fifo_cout_drain_out_V_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper497_U0_fifo_cout_drain_out_V_V_write_pass_1_q0 <= cout_drain_IO_L1_out_wrapper497_U0_fifo_cout_drain_out_V_V_write_pass_1_out;
  end
  assign cout_drain_IO_L1_out_wrapper497_U0_fifo_cout_drain_out_V_V_write_pass_1_in = cout_drain_IO_L1_out_wrapper497_U0_fifo_cout_drain_out_V_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper278_U0_fifo_w_out_V_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper278_U0_fifo_w_out_V_V_din_pass_1_q0 <= PE_wrapper278_U0_fifo_w_out_V_V_din_pass_1_out;
  end
  assign PE_wrapper278_U0_fifo_w_out_V_V_din_pass_1_in = PE_wrapper278_U0_fifo_w_out_V_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_10_9_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_10_9_V_V_full_n_pass_0_q0 <= fifo_w_PE_10_9_V_V_full_n_pass_0_out;
  end
  assign fifo_w_PE_10_9_V_V_full_n_pass_0_in = fifo_w_PE_10_9_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper278_U0_fifo_w_out_V_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper278_U0_fifo_w_out_V_V_write_pass_1_q0 <= PE_wrapper278_U0_fifo_w_out_V_V_write_pass_1_out;
  end
  assign PE_wrapper278_U0_fifo_w_out_V_V_write_pass_1_in = PE_wrapper278_U0_fifo_w_out_V_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_11_9_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_11_9_V_V_full_n_pass_0_q0 <= fifo_w_PE_11_9_V_V_full_n_pass_0_out;
  end
  assign fifo_w_PE_11_9_V_V_full_n_pass_0_in = fifo_w_PE_11_9_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper304_U0_fifo_cin_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper304_U0_fifo_cin_out_V_V_din_pass_0_q0 <= PE_wrapper304_U0_fifo_cin_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper304_U0_fifo_cin_out_V_V_din_pass_0_in = PE_wrapper304_U0_fifo_cin_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper304_U0_fifo_cin_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper304_U0_fifo_cin_out_V_V_write_pass_0_q0 <= PE_wrapper304_U0_fifo_cin_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper304_U0_fifo_cin_out_V_V_write_pass_0_in = PE_wrapper304_U0_fifo_cin_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_11_9_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_11_9_V_V_full_n_pass_0_q0 <= fifo_cin_PE_11_9_V_V_full_n_pass_0_out;
  end
  assign fifo_cin_PE_11_9_V_V_full_n_pass_0_in = fifo_cin_PE_11_9_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper267_U0_fifo_cin_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper267_U0_fifo_cin_out_V_V_din_pass_0_q0 <= PE_wrapper267_U0_fifo_cin_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper267_U0_fifo_cin_out_V_V_din_pass_0_in = PE_wrapper267_U0_fifo_cin_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper267_U0_fifo_cin_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper267_U0_fifo_cin_out_V_V_write_pass_0_q0 <= PE_wrapper267_U0_fifo_cin_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper267_U0_fifo_cin_out_V_V_write_pass_0_in = PE_wrapper267_U0_fifo_cin_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_PE_9_11_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_PE_9_11_V_full_n_pass_0_q0 <= fifo_cout_drain_PE_9_11_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_PE_9_11_V_full_n_pass_0_in = fifo_cout_drain_PE_9_11_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_cout_drain_IO_L1_out_9_13_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_cout_drain_IO_L1_out_9_13_V_V_full_n_pass_0_q0 <= fifo_cout_drain_cout_drain_IO_L1_out_9_13_V_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_cout_drain_IO_L1_out_9_13_V_V_full_n_pass_0_in = fifo_cout_drain_cout_drain_IO_L1_out_9_13_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_11_11_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_11_11_V_V_full_n_pass_0_q0 <= fifo_w_PE_11_11_V_V_full_n_pass_0_out;
  end
  assign fifo_w_PE_11_11_V_V_full_n_pass_0_in = fifo_w_PE_11_11_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_PE_10_11_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_PE_10_11_V_full_n_pass_0_q0 <= fifo_cout_drain_PE_10_11_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_PE_10_11_V_full_n_pass_0_in = fifo_cout_drain_PE_10_11_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_PE_10_10_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_PE_10_10_V_full_n_pass_0_q0 <= fifo_cout_drain_PE_10_10_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_PE_10_10_V_full_n_pass_0_in = fifo_cout_drain_PE_10_10_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_11_11_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_11_11_V_V_full_n_pass_0_q0 <= fifo_cin_PE_11_11_V_V_full_n_pass_0_out;
  end
  assign fifo_cin_PE_11_11_V_V_full_n_pass_0_in = fifo_cin_PE_11_11_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_12_9_V_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_12_9_V_V_full_n_pass_1_q0 <= fifo_w_PE_12_9_V_V_full_n_pass_1_out;
  end
  assign fifo_w_PE_12_9_V_V_full_n_pass_1_in = fifo_w_PE_12_9_V_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper291_U0_fifo_w_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper291_U0_fifo_w_out_V_V_din_pass_0_q0 <= PE_wrapper291_U0_fifo_w_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper291_U0_fifo_w_out_V_V_din_pass_0_in = PE_wrapper291_U0_fifo_w_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper291_U0_fifo_w_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper291_U0_fifo_w_out_V_V_write_pass_0_q0 <= PE_wrapper291_U0_fifo_w_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper291_U0_fifo_w_out_V_V_write_pass_0_in = PE_wrapper291_U0_fifo_w_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_9_9_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_9_9_V_V_full_n_pass_0_q0 <= fifo_cin_PE_9_9_V_V_full_n_pass_0_out;
  end
  assign fifo_cin_PE_9_9_V_V_full_n_pass_0_in = fifo_cin_PE_9_9_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_12_10_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_12_10_V_V_full_n_pass_0_q0 <= fifo_cin_PE_12_10_V_V_full_n_pass_0_out;
  end
  assign fifo_cin_PE_12_10_V_V_full_n_pass_0_in = fifo_cin_PE_12_10_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg [63:0] cout_drain_IO_L1_out_wrapper517_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper517_U0_fifo_cout_drain_out_V_V_din_pass_0_q0 <= cout_drain_IO_L1_out_wrapper517_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper517_U0_fifo_cout_drain_out_V_V_din_pass_0_in = cout_drain_IO_L1_out_wrapper517_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  cout_drain_IO_L1_out_wrapper517_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper517_U0_fifo_cout_drain_out_V_V_write_pass_0_q0 <= cout_drain_IO_L1_out_wrapper517_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper517_U0_fifo_cout_drain_out_V_V_write_pass_0_in = cout_drain_IO_L1_out_wrapper517_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_PE_9_10_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_PE_9_10_V_full_n_pass_0_q0 <= fifo_cout_drain_PE_9_10_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_PE_9_10_V_full_n_pass_0_in = fifo_cout_drain_PE_9_10_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_9_9_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_9_9_V_V_full_n_pass_0_q0 <= fifo_w_PE_9_9_V_V_full_n_pass_0_out;
  end
  assign fifo_w_PE_9_9_V_V_full_n_pass_0_in = fifo_w_PE_9_9_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_cout_drain_IO_L1_out_10_13_V_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_cout_drain_IO_L1_out_10_13_V_V_full_n_pass_1_q0 <= fifo_cout_drain_cout_drain_IO_L1_out_10_13_V_V_full_n_pass_1_out;
  end
  assign fifo_cout_drain_cout_drain_IO_L1_out_10_13_V_V_full_n_pass_1_in = fifo_cout_drain_cout_drain_IO_L1_out_10_13_V_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg [63:0] cout_drain_IO_L1_out_wrapper533_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper533_U0_fifo_cout_drain_out_V_V_din_pass_0_q0 <= cout_drain_IO_L1_out_wrapper533_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper533_U0_fifo_cout_drain_out_V_V_din_pass_0_in = cout_drain_IO_L1_out_wrapper533_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  cout_drain_IO_L1_out_wrapper533_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper533_U0_fifo_cout_drain_out_V_V_write_pass_0_q0 <= cout_drain_IO_L1_out_wrapper533_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper533_U0_fifo_cout_drain_out_V_V_write_pass_0_in = cout_drain_IO_L1_out_wrapper533_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper267_U0_fifo_w_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper267_U0_fifo_w_out_V_V_din_pass_0_q0 <= PE_wrapper267_U0_fifo_w_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper267_U0_fifo_w_out_V_V_din_pass_0_in = PE_wrapper267_U0_fifo_w_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper267_U0_fifo_w_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper267_U0_fifo_w_out_V_V_write_pass_0_q0 <= PE_wrapper267_U0_fifo_w_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper267_U0_fifo_w_out_V_V_write_pass_0_in = PE_wrapper267_U0_fifo_w_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper305_U0_fifo_cin_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper305_U0_fifo_cin_out_V_V_din_pass_0_q0 <= PE_wrapper305_U0_fifo_cin_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper305_U0_fifo_cin_out_V_V_din_pass_0_in = PE_wrapper305_U0_fifo_cin_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper305_U0_fifo_cin_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper305_U0_fifo_cin_out_V_V_write_pass_0_q0 <= PE_wrapper305_U0_fifo_cin_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper305_U0_fifo_cin_out_V_V_write_pass_0_in = PE_wrapper305_U0_fifo_cin_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_PE_11_10_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_PE_11_10_V_full_n_pass_0_q0 <= fifo_cout_drain_PE_11_10_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_PE_11_10_V_full_n_pass_0_in = fifo_cout_drain_PE_11_10_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg [63:0] cout_drain_IO_L1_out_wrapper548_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper548_U0_fifo_cout_drain_out_V_V_din_pass_0_q0 <= cout_drain_IO_L1_out_wrapper548_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper548_U0_fifo_cout_drain_out_V_V_din_pass_0_in = cout_drain_IO_L1_out_wrapper548_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  cout_drain_IO_L1_out_wrapper548_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper548_U0_fifo_cout_drain_out_V_V_write_pass_0_q0 <= cout_drain_IO_L1_out_wrapper548_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper548_U0_fifo_cout_drain_out_V_V_write_pass_0_in = cout_drain_IO_L1_out_wrapper548_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_PE_10_9_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_PE_10_9_V_full_n_pass_0_q0 <= fifo_cout_drain_PE_10_9_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_PE_10_9_V_full_n_pass_0_in = fifo_cout_drain_PE_10_9_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper303_U0_fifo_cin_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper303_U0_fifo_cin_out_V_V_din_pass_0_q0 <= PE_wrapper303_U0_fifo_cin_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper303_U0_fifo_cin_out_V_V_din_pass_0_in = PE_wrapper303_U0_fifo_cin_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper303_U0_fifo_cin_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper303_U0_fifo_cin_out_V_V_write_pass_0_q0 <= PE_wrapper303_U0_fifo_cin_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper303_U0_fifo_cin_out_V_V_write_pass_0_in = PE_wrapper303_U0_fifo_cin_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_cout_drain_IO_L1_out_11_13_V_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_cout_drain_IO_L1_out_11_13_V_V_full_n_pass_1_q0 <= fifo_cout_drain_cout_drain_IO_L1_out_11_13_V_V_full_n_pass_1_out;
  end
  assign fifo_cout_drain_cout_drain_IO_L1_out_11_13_V_V_full_n_pass_1_in = fifo_cout_drain_cout_drain_IO_L1_out_11_13_V_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg  ap_done_Boundary_X2Y12_To_X4Y12_q0;
  always @ (posedge ap_clk) begin
    ap_done_Boundary_X2Y12_To_X4Y12_q0 <= ap_done_Boundary_X2Y12_To_X4Y12_out;
  end
  assign ap_done_Boundary_X2Y12_To_X4Y12_in = ap_done_Boundary_X2Y12_To_X4Y12_q0;
  (* dont_touch = "yes" *) reg  ap_start_Boundary_X2Y14_To_X4Y14_q0;
  always @ (posedge ap_clk) begin
    ap_start_Boundary_X2Y14_To_X4Y14_q0 <= ap_start_Boundary_X2Y14_To_X4Y14_out;
  end
  assign ap_start_Boundary_X2Y14_To_X4Y14_in = ap_start_Boundary_X2Y14_To_X4Y14_q0;
  (* dont_touch = "yes" *) reg  ap_rst_n_Boundary_X2Y14_To_X4Y14_q0;
  always @ (posedge ap_clk) begin
    ap_rst_n_Boundary_X2Y14_To_X4Y14_q0 <= ap_rst_n_Boundary_X2Y14_To_X4Y14_out;
  end
  assign ap_rst_n_Boundary_X2Y14_To_X4Y14_in = ap_rst_n_Boundary_X2Y14_To_X4Y14_q0;
  (* dont_touch = "yes" *) reg [63:0] cout_drain_IO_L1_out_wrapper529_U0_fifo_cout_drain_out_V_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper529_U0_fifo_cout_drain_out_V_V_din_pass_1_q0 <= cout_drain_IO_L1_out_wrapper529_U0_fifo_cout_drain_out_V_V_din_pass_1_out;
  end
  assign cout_drain_IO_L1_out_wrapper529_U0_fifo_cout_drain_out_V_V_din_pass_1_in = cout_drain_IO_L1_out_wrapper529_U0_fifo_cout_drain_out_V_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_cout_drain_IO_L1_out_10_13_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_cout_drain_IO_L1_out_10_13_V_V_full_n_pass_0_q0 <= fifo_cout_drain_cout_drain_IO_L1_out_10_13_V_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_cout_drain_IO_L1_out_10_13_V_V_full_n_pass_0_in = fifo_cout_drain_cout_drain_IO_L1_out_10_13_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  cout_drain_IO_L1_out_wrapper529_U0_fifo_cout_drain_out_V_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper529_U0_fifo_cout_drain_out_V_V_write_pass_1_q0 <= cout_drain_IO_L1_out_wrapper529_U0_fifo_cout_drain_out_V_V_write_pass_1_out;
  end
  assign cout_drain_IO_L1_out_wrapper529_U0_fifo_cout_drain_out_V_V_write_pass_1_in = cout_drain_IO_L1_out_wrapper529_U0_fifo_cout_drain_out_V_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [63:0] cout_drain_IO_L1_out_wrapper544_U0_fifo_cout_drain_out_V_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper544_U0_fifo_cout_drain_out_V_V_din_pass_1_q0 <= cout_drain_IO_L1_out_wrapper544_U0_fifo_cout_drain_out_V_V_din_pass_1_out;
  end
  assign cout_drain_IO_L1_out_wrapper544_U0_fifo_cout_drain_out_V_V_din_pass_1_in = cout_drain_IO_L1_out_wrapper544_U0_fifo_cout_drain_out_V_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_cout_drain_IO_L1_out_11_13_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_cout_drain_IO_L1_out_11_13_V_V_full_n_pass_0_q0 <= fifo_cout_drain_cout_drain_IO_L1_out_11_13_V_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_cout_drain_IO_L1_out_11_13_V_V_full_n_pass_0_in = fifo_cout_drain_cout_drain_IO_L1_out_11_13_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  cout_drain_IO_L1_out_wrapper544_U0_fifo_cout_drain_out_V_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper544_U0_fifo_cout_drain_out_V_V_write_pass_1_q0 <= cout_drain_IO_L1_out_wrapper544_U0_fifo_cout_drain_out_V_V_write_pass_1_out;
  end
  assign cout_drain_IO_L1_out_wrapper544_U0_fifo_cout_drain_out_V_V_write_pass_1_in = cout_drain_IO_L1_out_wrapper544_U0_fifo_cout_drain_out_V_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper279_U0_fifo_cin_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper279_U0_fifo_cin_out_V_V_din_pass_0_q0 <= PE_wrapper279_U0_fifo_cin_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper279_U0_fifo_cin_out_V_V_din_pass_0_in = PE_wrapper279_U0_fifo_cin_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper279_U0_fifo_cin_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper279_U0_fifo_cin_out_V_V_write_pass_0_q0 <= PE_wrapper279_U0_fifo_cin_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper279_U0_fifo_cin_out_V_V_write_pass_0_in = PE_wrapper279_U0_fifo_cin_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [31:0] PE_wrapper269_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper269_U0_fifo_cout_drain_out_V_din_pass_0_q0 <= PE_wrapper269_U0_fifo_cout_drain_out_V_din_pass_0_out;
  end
  assign PE_wrapper269_U0_fifo_cout_drain_out_V_din_pass_0_in = PE_wrapper269_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper269_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper269_U0_fifo_cout_drain_out_V_write_pass_0_q0 <= PE_wrapper269_U0_fifo_cout_drain_out_V_write_pass_0_out;
  end
  assign PE_wrapper269_U0_fifo_cout_drain_out_V_write_pass_0_in = PE_wrapper269_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_10_9_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_10_9_V_V_full_n_pass_0_q0 <= fifo_cin_PE_10_9_V_V_full_n_pass_0_out;
  end
  assign fifo_cin_PE_10_9_V_V_full_n_pass_0_in = fifo_cin_PE_10_9_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper292_U0_fifo_w_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper292_U0_fifo_w_out_V_V_din_pass_0_q0 <= PE_wrapper292_U0_fifo_w_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper292_U0_fifo_w_out_V_V_din_pass_0_in = PE_wrapper292_U0_fifo_w_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper292_U0_fifo_w_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper292_U0_fifo_w_out_V_V_write_pass_0_q0 <= PE_wrapper292_U0_fifo_w_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper292_U0_fifo_w_out_V_V_write_pass_0_in = PE_wrapper292_U0_fifo_w_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [31:0] PE_wrapper281_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper281_U0_fifo_cout_drain_out_V_din_pass_0_q0 <= PE_wrapper281_U0_fifo_cout_drain_out_V_din_pass_0_out;
  end
  assign PE_wrapper281_U0_fifo_cout_drain_out_V_din_pass_0_in = PE_wrapper281_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper281_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper281_U0_fifo_cout_drain_out_V_write_pass_0_q0 <= PE_wrapper281_U0_fifo_cout_drain_out_V_write_pass_0_out;
  end
  assign PE_wrapper281_U0_fifo_cout_drain_out_V_write_pass_0_in = PE_wrapper281_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [31:0] PE_wrapper280_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper280_U0_fifo_cout_drain_out_V_din_pass_0_q0 <= PE_wrapper280_U0_fifo_cout_drain_out_V_din_pass_0_out;
  end
  assign PE_wrapper280_U0_fifo_cout_drain_out_V_din_pass_0_in = PE_wrapper280_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper280_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper280_U0_fifo_cout_drain_out_V_write_pass_0_q0 <= PE_wrapper280_U0_fifo_cout_drain_out_V_write_pass_0_out;
  end
  assign PE_wrapper280_U0_fifo_cout_drain_out_V_write_pass_0_in = PE_wrapper280_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_10_9_V_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_10_9_V_V_full_n_pass_1_q0 <= fifo_w_PE_10_9_V_V_full_n_pass_1_out;
  end
  assign fifo_w_PE_10_9_V_V_full_n_pass_1_in = fifo_w_PE_10_9_V_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper281_U0_fifo_cin_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper281_U0_fifo_cin_out_V_V_din_pass_0_q0 <= PE_wrapper281_U0_fifo_cin_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper281_U0_fifo_cin_out_V_V_din_pass_0_in = PE_wrapper281_U0_fifo_cin_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper281_U0_fifo_cin_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper281_U0_fifo_cin_out_V_V_write_pass_0_q0 <= PE_wrapper281_U0_fifo_cin_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper281_U0_fifo_cin_out_V_V_write_pass_0_in = PE_wrapper281_U0_fifo_cin_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_9_10_V_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_9_10_V_V_full_n_pass_1_q0 <= fifo_cin_PE_9_10_V_V_full_n_pass_1_out;
  end
  assign fifo_cin_PE_9_10_V_V_full_n_pass_1_in = fifo_cin_PE_9_10_V_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_11_10_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_11_10_V_V_full_n_pass_0_q0 <= fifo_w_PE_11_10_V_V_full_n_pass_0_out;
  end
  assign fifo_w_PE_11_10_V_V_full_n_pass_0_in = fifo_w_PE_11_10_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper292_U0_fifo_cin_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper292_U0_fifo_cin_out_V_V_din_pass_0_q0 <= PE_wrapper292_U0_fifo_cin_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper292_U0_fifo_cin_out_V_V_din_pass_0_in = PE_wrapper292_U0_fifo_cin_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper292_U0_fifo_cin_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper292_U0_fifo_cin_out_V_V_write_pass_0_q0 <= PE_wrapper292_U0_fifo_cin_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper292_U0_fifo_cin_out_V_V_write_pass_0_in = PE_wrapper292_U0_fifo_cin_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [31:0] PE_wrapper268_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper268_U0_fifo_cout_drain_out_V_din_pass_0_q0 <= PE_wrapper268_U0_fifo_cout_drain_out_V_din_pass_0_out;
  end
  assign PE_wrapper268_U0_fifo_cout_drain_out_V_din_pass_0_in = PE_wrapper268_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper268_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper268_U0_fifo_cout_drain_out_V_write_pass_0_q0 <= PE_wrapper268_U0_fifo_cout_drain_out_V_write_pass_0_out;
  end
  assign PE_wrapper268_U0_fifo_cout_drain_out_V_write_pass_0_in = PE_wrapper268_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_9_11_V_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_9_11_V_V_full_n_pass_1_q0 <= fifo_cin_PE_9_11_V_V_full_n_pass_1_out;
  end
  assign fifo_cin_PE_9_11_V_V_full_n_pass_1_in = fifo_cin_PE_9_11_V_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_9_10_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_9_10_V_V_full_n_pass_0_q0 <= fifo_w_PE_9_10_V_V_full_n_pass_0_out;
  end
  assign fifo_w_PE_9_10_V_V_full_n_pass_0_in = fifo_w_PE_9_10_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg [31:0] PE_wrapper292_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper292_U0_fifo_cout_drain_out_V_din_pass_0_q0 <= PE_wrapper292_U0_fifo_cout_drain_out_V_din_pass_0_out;
  end
  assign PE_wrapper292_U0_fifo_cout_drain_out_V_din_pass_0_in = PE_wrapper292_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper292_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper292_U0_fifo_cout_drain_out_V_write_pass_0_q0 <= PE_wrapper292_U0_fifo_cout_drain_out_V_write_pass_0_out;
  end
  assign PE_wrapper292_U0_fifo_cout_drain_out_V_write_pass_0_in = PE_wrapper292_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [31:0] PE_wrapper279_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper279_U0_fifo_cout_drain_out_V_din_pass_0_q0 <= PE_wrapper279_U0_fifo_cout_drain_out_V_din_pass_0_out;
  end
  assign PE_wrapper279_U0_fifo_cout_drain_out_V_din_pass_0_in = PE_wrapper279_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper279_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper279_U0_fifo_cout_drain_out_V_write_pass_0_q0 <= PE_wrapper279_U0_fifo_cout_drain_out_V_write_pass_0_out;
  end
  assign PE_wrapper279_U0_fifo_cout_drain_out_V_write_pass_0_in = PE_wrapper279_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  ap_done_Boundary_X2Y14_To_X4Y14_q0;
  always @ (posedge ap_clk) begin
    ap_done_Boundary_X2Y14_To_X4Y14_q0 <= ap_done_Boundary_X2Y14_To_X4Y14_out;
  end
  assign ap_done_Boundary_X2Y14_To_X4Y14_in = ap_done_Boundary_X2Y14_To_X4Y14_q0;
  (* dont_touch = "yes" *) reg [255:0] w_IO_L2_in140_U0_fifo_w_out_V_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    w_IO_L2_in140_U0_fifo_w_out_V_V_din_pass_1_q0 <= w_IO_L2_in140_U0_fifo_w_out_V_V_din_pass_1_out;
  end
  assign w_IO_L2_in140_U0_fifo_w_out_V_V_din_pass_1_in = w_IO_L2_in140_U0_fifo_w_out_V_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_w_w_IO_L2_in_6_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_w_IO_L2_in_6_V_V_full_n_pass_0_q0 <= fifo_w_w_IO_L2_in_6_V_V_full_n_pass_0_out;
  end
  assign fifo_w_w_IO_L2_in_6_V_V_full_n_pass_0_in = fifo_w_w_IO_L2_in_6_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  w_IO_L2_in140_U0_fifo_w_out_V_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    w_IO_L2_in140_U0_fifo_w_out_V_V_write_pass_1_q0 <= w_IO_L2_in140_U0_fifo_w_out_V_V_write_pass_1_out;
  end
  assign w_IO_L2_in140_U0_fifo_w_out_V_V_write_pass_1_in = w_IO_L2_in140_U0_fifo_w_out_V_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper210_U0_fifo_cin_out_V_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper210_U0_fifo_cin_out_V_V_din_pass_1_q0 <= PE_wrapper210_U0_fifo_cin_out_V_V_din_pass_1_out;
  end
  assign PE_wrapper210_U0_fifo_cin_out_V_V_din_pass_1_in = PE_wrapper210_U0_fifo_cin_out_V_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_6_0_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_6_0_V_V_full_n_pass_0_q0 <= fifo_cin_PE_6_0_V_V_full_n_pass_0_out;
  end
  assign fifo_cin_PE_6_0_V_V_full_n_pass_0_in = fifo_cin_PE_6_0_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper210_U0_fifo_cin_out_V_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper210_U0_fifo_cin_out_V_V_write_pass_1_q0 <= PE_wrapper210_U0_fifo_cin_out_V_V_write_pass_1_out;
  end
  assign PE_wrapper210_U0_fifo_cin_out_V_V_write_pass_1_in = PE_wrapper210_U0_fifo_cin_out_V_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [255:0] w_IO_L2_in138_U0_fifo_w_local_out_V_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    w_IO_L2_in138_U0_fifo_w_local_out_V_V_din_pass_1_q0 <= w_IO_L2_in138_U0_fifo_w_local_out_V_V_din_pass_1_out;
  end
  assign w_IO_L2_in138_U0_fifo_w_local_out_V_V_din_pass_1_in = w_IO_L2_in138_U0_fifo_w_local_out_V_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_3_0_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_3_0_V_V_full_n_pass_0_q0 <= fifo_w_PE_3_0_V_V_full_n_pass_0_out;
  end
  assign fifo_w_PE_3_0_V_V_full_n_pass_0_in = fifo_w_PE_3_0_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  w_IO_L2_in138_U0_fifo_w_local_out_V_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    w_IO_L2_in138_U0_fifo_w_local_out_V_V_write_pass_1_q0 <= w_IO_L2_in138_U0_fifo_w_local_out_V_V_write_pass_1_out;
  end
  assign w_IO_L2_in138_U0_fifo_w_local_out_V_V_write_pass_1_in = w_IO_L2_in138_U0_fifo_w_local_out_V_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [63:0] cout_drain_IO_L1_out_wrapper378_U0_fifo_cout_drain_out_V_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper378_U0_fifo_cout_drain_out_V_V_din_pass_1_q0 <= cout_drain_IO_L1_out_wrapper378_U0_fifo_cout_drain_out_V_V_din_pass_1_out;
  end
  assign cout_drain_IO_L1_out_wrapper378_U0_fifo_cout_drain_out_V_V_din_pass_1_in = cout_drain_IO_L1_out_wrapper378_U0_fifo_cout_drain_out_V_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_cout_drain_IO_L1_out_0_4_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_cout_drain_IO_L1_out_0_4_V_V_full_n_pass_0_q0 <= fifo_cout_drain_cout_drain_IO_L1_out_0_4_V_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_cout_drain_IO_L1_out_0_4_V_V_full_n_pass_0_in = fifo_cout_drain_cout_drain_IO_L1_out_0_4_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  cout_drain_IO_L1_out_wrapper378_U0_fifo_cout_drain_out_V_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper378_U0_fifo_cout_drain_out_V_V_write_pass_1_q0 <= cout_drain_IO_L1_out_wrapper378_U0_fifo_cout_drain_out_V_V_write_pass_1_out;
  end
  assign cout_drain_IO_L1_out_wrapper378_U0_fifo_cout_drain_out_V_V_write_pass_1_in = cout_drain_IO_L1_out_wrapper378_U0_fifo_cout_drain_out_V_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper201_U0_fifo_w_out_V_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper201_U0_fifo_w_out_V_V_din_pass_1_q0 <= PE_wrapper201_U0_fifo_w_out_V_V_din_pass_1_out;
  end
  assign PE_wrapper201_U0_fifo_w_out_V_V_din_pass_1_in = PE_wrapper201_U0_fifo_w_out_V_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_4_4_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_4_4_V_V_full_n_pass_0_q0 <= fifo_w_PE_4_4_V_V_full_n_pass_0_out;
  end
  assign fifo_w_PE_4_4_V_V_full_n_pass_0_in = fifo_w_PE_4_4_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper201_U0_fifo_w_out_V_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper201_U0_fifo_w_out_V_V_write_pass_1_q0 <= PE_wrapper201_U0_fifo_w_out_V_V_write_pass_1_out;
  end
  assign PE_wrapper201_U0_fifo_w_out_V_V_write_pass_1_in = PE_wrapper201_U0_fifo_w_out_V_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper213_U0_fifo_w_out_V_V_din_pass_2_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper213_U0_fifo_w_out_V_V_din_pass_2_q0 <= PE_wrapper213_U0_fifo_w_out_V_V_din_pass_2_out;
  end
  assign PE_wrapper213_U0_fifo_w_out_V_V_din_pass_2_in = PE_wrapper213_U0_fifo_w_out_V_V_din_pass_2_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_5_4_V_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_5_4_V_V_full_n_pass_1_q0 <= fifo_w_PE_5_4_V_V_full_n_pass_1_out;
  end
  assign fifo_w_PE_5_4_V_V_full_n_pass_1_in = fifo_w_PE_5_4_V_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper213_U0_fifo_w_out_V_V_write_pass_2_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper213_U0_fifo_w_out_V_V_write_pass_2_q0 <= PE_wrapper213_U0_fifo_w_out_V_V_write_pass_2_out;
  end
  assign PE_wrapper213_U0_fifo_w_out_V_V_write_pass_2_in = PE_wrapper213_U0_fifo_w_out_V_V_write_pass_2_q0;
  (* dont_touch = "yes" *) reg [63:0] kernel0_entry12_U0_w_V_out_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    kernel0_entry12_U0_w_V_out_din_pass_1_q0 <= kernel0_entry12_U0_w_V_out_din_pass_1_out;
  end
  assign kernel0_entry12_U0_w_V_out_din_pass_1_in = kernel0_entry12_U0_w_V_out_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  w_V_c_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    w_V_c_full_n_pass_0_q0 <= w_V_c_full_n_pass_0_out;
  end
  assign w_V_c_full_n_pass_0_in = w_V_c_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  kernel0_entry12_U0_w_V_out_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    kernel0_entry12_U0_w_V_out_write_pass_1_q0 <= kernel0_entry12_U0_w_V_out_write_pass_1_out;
  end
  assign kernel0_entry12_U0_w_V_out_write_pass_1_in = kernel0_entry12_U0_w_V_out_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [63:0] kernel0_entry12_U0_cout_V_out_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    kernel0_entry12_U0_cout_V_out_din_pass_1_q0 <= kernel0_entry12_U0_cout_V_out_din_pass_1_out;
  end
  assign kernel0_entry12_U0_cout_V_out_din_pass_1_in = kernel0_entry12_U0_cout_V_out_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  cout_V_c_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_V_c_full_n_pass_0_q0 <= cout_V_c_full_n_pass_0_out;
  end
  assign cout_V_c_full_n_pass_0_in = cout_V_c_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  kernel0_entry12_U0_cout_V_out_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    kernel0_entry12_U0_cout_V_out_write_pass_1_q0 <= kernel0_entry12_U0_cout_V_out_write_pass_1_out;
  end
  assign kernel0_entry12_U0_cout_V_out_write_pass_1_in = kernel0_entry12_U0_cout_V_out_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper165_U0_fifo_w_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper165_U0_fifo_w_out_V_V_din_pass_0_q0 <= PE_wrapper165_U0_fifo_w_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper165_U0_fifo_w_out_V_V_din_pass_0_in = PE_wrapper165_U0_fifo_w_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper165_U0_fifo_w_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper165_U0_fifo_w_out_V_V_write_pass_0_q0 <= PE_wrapper165_U0_fifo_w_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper165_U0_fifo_w_out_V_V_write_pass_0_in = PE_wrapper165_U0_fifo_w_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] cin_IO_L2_in127_U0_fifo_cin_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    cin_IO_L2_in127_U0_fifo_cin_out_V_V_din_pass_0_q0 <= cin_IO_L2_in127_U0_fifo_cin_out_V_V_din_pass_0_out;
  end
  assign cin_IO_L2_in127_U0_fifo_cin_out_V_V_din_pass_0_in = cin_IO_L2_in127_U0_fifo_cin_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  cin_IO_L2_in127_U0_fifo_cin_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    cin_IO_L2_in127_U0_fifo_cin_out_V_V_write_pass_0_q0 <= cin_IO_L2_in127_U0_fifo_cin_out_V_V_write_pass_0_out;
  end
  assign cin_IO_L2_in127_U0_fifo_cin_out_V_V_write_pass_0_in = cin_IO_L2_in127_U0_fifo_cin_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_1_2_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_1_2_V_V_full_n_pass_0_q0 <= fifo_w_PE_1_2_V_V_full_n_pass_0_out;
  end
  assign fifo_w_PE_1_2_V_V_full_n_pass_0_in = fifo_w_PE_1_2_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_3_3_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_3_3_V_V_full_n_pass_0_q0 <= fifo_w_PE_3_3_V_V_full_n_pass_0_out;
  end
  assign fifo_w_PE_3_3_V_V_full_n_pass_0_in = fifo_w_PE_3_3_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] w_IO_L2_in136_U0_fifo_w_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    w_IO_L2_in136_U0_fifo_w_out_V_V_din_pass_0_q0 <= w_IO_L2_in136_U0_fifo_w_out_V_V_din_pass_0_out;
  end
  assign w_IO_L2_in136_U0_fifo_w_out_V_V_din_pass_0_in = w_IO_L2_in136_U0_fifo_w_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  w_IO_L2_in136_U0_fifo_w_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    w_IO_L2_in136_U0_fifo_w_out_V_V_write_pass_0_q0 <= w_IO_L2_in136_U0_fifo_w_out_V_V_write_pass_0_out;
  end
  assign w_IO_L2_in136_U0_fifo_w_out_V_V_write_pass_0_in = w_IO_L2_in136_U0_fifo_w_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper153_U0_fifo_w_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper153_U0_fifo_w_out_V_V_din_pass_0_q0 <= PE_wrapper153_U0_fifo_w_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper153_U0_fifo_w_out_V_V_din_pass_0_in = PE_wrapper153_U0_fifo_w_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper153_U0_fifo_w_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper153_U0_fifo_w_out_V_V_write_pass_0_q0 <= PE_wrapper153_U0_fifo_w_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper153_U0_fifo_w_out_V_V_write_pass_0_in = PE_wrapper153_U0_fifo_w_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper177_U0_fifo_w_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper177_U0_fifo_w_out_V_V_din_pass_0_q0 <= PE_wrapper177_U0_fifo_w_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper177_U0_fifo_w_out_V_V_din_pass_0_in = PE_wrapper177_U0_fifo_w_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper177_U0_fifo_w_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper177_U0_fifo_w_out_V_V_write_pass_0_q0 <= PE_wrapper177_U0_fifo_w_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper177_U0_fifo_w_out_V_V_write_pass_0_in = PE_wrapper177_U0_fifo_w_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_0_2_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_0_2_V_V_full_n_pass_0_q0 <= fifo_w_PE_0_2_V_V_full_n_pass_0_out;
  end
  assign fifo_w_PE_0_2_V_V_full_n_pass_0_in = fifo_w_PE_0_2_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg [31:0] PE_wrapper165_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper165_U0_fifo_cout_drain_out_V_din_pass_0_q0 <= PE_wrapper165_U0_fifo_cout_drain_out_V_din_pass_0_out;
  end
  assign PE_wrapper165_U0_fifo_cout_drain_out_V_din_pass_0_in = PE_wrapper165_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper165_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper165_U0_fifo_cout_drain_out_V_write_pass_0_q0 <= PE_wrapper165_U0_fifo_cout_drain_out_V_write_pass_0_out;
  end
  assign PE_wrapper165_U0_fifo_cout_drain_out_V_write_pass_0_in = PE_wrapper165_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_1_0_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_1_0_V_V_full_n_pass_0_q0 <= fifo_cin_PE_1_0_V_V_full_n_pass_0_out;
  end
  assign fifo_cin_PE_1_0_V_V_full_n_pass_0_in = fifo_cin_PE_1_0_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg [31:0] PE_wrapper153_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper153_U0_fifo_cout_drain_out_V_din_pass_0_q0 <= PE_wrapper153_U0_fifo_cout_drain_out_V_din_pass_0_out;
  end
  assign PE_wrapper153_U0_fifo_cout_drain_out_V_din_pass_0_in = PE_wrapper153_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper153_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper153_U0_fifo_cout_drain_out_V_write_pass_0_q0 <= PE_wrapper153_U0_fifo_cout_drain_out_V_write_pass_0_out;
  end
  assign PE_wrapper153_U0_fifo_cout_drain_out_V_write_pass_0_in = PE_wrapper153_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [31:0] PE_wrapper177_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper177_U0_fifo_cout_drain_out_V_din_pass_0_q0 <= PE_wrapper177_U0_fifo_cout_drain_out_V_din_pass_0_out;
  end
  assign PE_wrapper177_U0_fifo_cout_drain_out_V_din_pass_0_in = PE_wrapper177_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper177_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper177_U0_fifo_cout_drain_out_V_write_pass_0_q0 <= PE_wrapper177_U0_fifo_cout_drain_out_V_write_pass_0_out;
  end
  assign PE_wrapper177_U0_fifo_cout_drain_out_V_write_pass_0_in = PE_wrapper177_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [31:0] PE_wrapper164_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper164_U0_fifo_cout_drain_out_V_din_pass_0_q0 <= PE_wrapper164_U0_fifo_cout_drain_out_V_din_pass_0_out;
  end
  assign PE_wrapper164_U0_fifo_cout_drain_out_V_din_pass_0_in = PE_wrapper164_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper164_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper164_U0_fifo_cout_drain_out_V_write_pass_0_q0 <= PE_wrapper164_U0_fifo_cout_drain_out_V_write_pass_0_out;
  end
  assign PE_wrapper164_U0_fifo_cout_drain_out_V_write_pass_0_in = PE_wrapper164_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [31:0] PE_wrapper189_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper189_U0_fifo_cout_drain_out_V_din_pass_0_q0 <= PE_wrapper189_U0_fifo_cout_drain_out_V_din_pass_0_out;
  end
  assign PE_wrapper189_U0_fifo_cout_drain_out_V_din_pass_0_in = PE_wrapper189_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper189_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper189_U0_fifo_cout_drain_out_V_write_pass_0_q0 <= PE_wrapper189_U0_fifo_cout_drain_out_V_write_pass_0_out;
  end
  assign PE_wrapper189_U0_fifo_cout_drain_out_V_write_pass_0_in = PE_wrapper189_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper162_U0_fifo_cin_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper162_U0_fifo_cin_out_V_V_din_pass_0_q0 <= PE_wrapper162_U0_fifo_cin_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper162_U0_fifo_cin_out_V_V_din_pass_0_in = PE_wrapper162_U0_fifo_cin_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper162_U0_fifo_cin_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper162_U0_fifo_cin_out_V_V_write_pass_0_q0 <= PE_wrapper162_U0_fifo_cin_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper162_U0_fifo_cin_out_V_V_write_pass_0_in = PE_wrapper162_U0_fifo_cin_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_w_w_IO_L3_in_serialize_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_w_IO_L3_in_serialize_V_V_full_n_pass_0_q0 <= fifo_w_w_IO_L3_in_serialize_V_V_full_n_pass_0_out;
  end
  assign fifo_w_w_IO_L3_in_serialize_V_V_full_n_pass_0_in = fifo_w_w_IO_L3_in_serialize_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_cin_IO_L2_in_2_V_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_cin_IO_L2_in_2_V_V_full_n_pass_1_q0 <= fifo_cin_cin_IO_L2_in_2_V_V_full_n_pass_1_out;
  end
  assign fifo_cin_cin_IO_L2_in_2_V_V_full_n_pass_1_in = fifo_cin_cin_IO_L2_in_2_V_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg [31:0] PE_wrapper152_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper152_U0_fifo_cout_drain_out_V_din_pass_0_q0 <= PE_wrapper152_U0_fifo_cout_drain_out_V_din_pass_0_out;
  end
  assign PE_wrapper152_U0_fifo_cout_drain_out_V_din_pass_0_in = PE_wrapper152_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper152_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper152_U0_fifo_cout_drain_out_V_write_pass_0_q0 <= PE_wrapper152_U0_fifo_cout_drain_out_V_write_pass_0_out;
  end
  assign PE_wrapper152_U0_fifo_cout_drain_out_V_write_pass_0_in = PE_wrapper152_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper189_U0_fifo_w_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper189_U0_fifo_w_out_V_V_din_pass_0_q0 <= PE_wrapper189_U0_fifo_w_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper189_U0_fifo_w_out_V_V_din_pass_0_in = PE_wrapper189_U0_fifo_w_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper189_U0_fifo_w_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper189_U0_fifo_w_out_V_V_write_pass_0_q0 <= PE_wrapper189_U0_fifo_w_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper189_U0_fifo_w_out_V_V_write_pass_0_in = PE_wrapper189_U0_fifo_w_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_2_2_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_2_2_V_V_full_n_pass_0_q0 <= fifo_w_PE_2_2_V_V_full_n_pass_0_out;
  end
  assign fifo_w_PE_2_2_V_V_full_n_pass_0_in = fifo_w_PE_2_2_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper162_U0_fifo_w_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper162_U0_fifo_w_out_V_V_din_pass_0_q0 <= PE_wrapper162_U0_fifo_w_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper162_U0_fifo_w_out_V_V_din_pass_0_in = PE_wrapper162_U0_fifo_w_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper162_U0_fifo_w_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper162_U0_fifo_w_out_V_V_write_pass_0_q0 <= PE_wrapper162_U0_fifo_w_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper162_U0_fifo_w_out_V_V_write_pass_0_in = PE_wrapper162_U0_fifo_w_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper189_U0_fifo_cin_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper189_U0_fifo_cin_out_V_V_din_pass_0_q0 <= PE_wrapper189_U0_fifo_cin_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper189_U0_fifo_cin_out_V_V_din_pass_0_in = PE_wrapper189_U0_fifo_cin_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper189_U0_fifo_cin_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper189_U0_fifo_cin_out_V_V_write_pass_0_q0 <= PE_wrapper189_U0_fifo_cin_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper189_U0_fifo_cin_out_V_V_write_pass_0_in = PE_wrapper189_U0_fifo_cin_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [31:0] PE_wrapper176_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper176_U0_fifo_cout_drain_out_V_din_pass_0_q0 <= PE_wrapper176_U0_fifo_cout_drain_out_V_din_pass_0_out;
  end
  assign PE_wrapper176_U0_fifo_cout_drain_out_V_din_pass_0_in = PE_wrapper176_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper176_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper176_U0_fifo_cout_drain_out_V_write_pass_0_q0 <= PE_wrapper176_U0_fifo_cout_drain_out_V_write_pass_0_out;
  end
  assign PE_wrapper176_U0_fifo_cout_drain_out_V_write_pass_0_in = PE_wrapper176_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper176_U0_fifo_cin_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper176_U0_fifo_cin_out_V_V_din_pass_0_q0 <= PE_wrapper176_U0_fifo_cin_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper176_U0_fifo_cin_out_V_V_din_pass_0_in = PE_wrapper176_U0_fifo_cin_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper176_U0_fifo_cin_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper176_U0_fifo_cin_out_V_V_write_pass_0_q0 <= PE_wrapper176_U0_fifo_cin_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper176_U0_fifo_cin_out_V_V_write_pass_0_in = PE_wrapper176_U0_fifo_cin_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [31:0] PE_wrapper162_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper162_U0_fifo_cout_drain_out_V_din_pass_0_q0 <= PE_wrapper162_U0_fifo_cout_drain_out_V_din_pass_0_out;
  end
  assign PE_wrapper162_U0_fifo_cout_drain_out_V_din_pass_0_in = PE_wrapper162_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper162_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper162_U0_fifo_cout_drain_out_V_write_pass_0_q0 <= PE_wrapper162_U0_fifo_cout_drain_out_V_write_pass_0_out;
  end
  assign PE_wrapper162_U0_fifo_cout_drain_out_V_write_pass_0_in = PE_wrapper162_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] w_IO_L2_in135_U0_fifo_w_local_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    w_IO_L2_in135_U0_fifo_w_local_out_V_V_din_pass_0_q0 <= w_IO_L2_in135_U0_fifo_w_local_out_V_V_din_pass_0_out;
  end
  assign w_IO_L2_in135_U0_fifo_w_local_out_V_V_din_pass_0_in = w_IO_L2_in135_U0_fifo_w_local_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  w_IO_L2_in135_U0_fifo_w_local_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    w_IO_L2_in135_U0_fifo_w_local_out_V_V_write_pass_0_q0 <= w_IO_L2_in135_U0_fifo_w_local_out_V_V_write_pass_0_out;
  end
  assign w_IO_L2_in135_U0_fifo_w_local_out_V_V_write_pass_0_in = w_IO_L2_in135_U0_fifo_w_local_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  ap_done_Boundary_X4Y2_To_X6Y2_q0;
  always @ (posedge ap_clk) begin
    ap_done_Boundary_X4Y2_To_X6Y2_q0 <= ap_done_Boundary_X4Y2_To_X6Y2_out;
  end
  assign ap_done_Boundary_X4Y2_To_X6Y2_in = ap_done_Boundary_X4Y2_To_X6Y2_q0;
  (* dont_touch = "yes" *) reg  ap_start_Boundary_X4Y4_To_X6Y4_q0;
  always @ (posedge ap_clk) begin
    ap_start_Boundary_X4Y4_To_X6Y4_q0 <= ap_start_Boundary_X4Y4_To_X6Y4_out;
  end
  assign ap_start_Boundary_X4Y4_To_X6Y4_in = ap_start_Boundary_X4Y4_To_X6Y4_q0;
  (* dont_touch = "yes" *) reg  ap_rst_n_Boundary_X4Y4_To_X6Y4_q0;
  always @ (posedge ap_clk) begin
    ap_rst_n_Boundary_X4Y4_To_X6Y4_q0 <= ap_rst_n_Boundary_X4Y4_To_X6Y4_out;
  end
  assign ap_rst_n_Boundary_X4Y4_To_X6Y4_in = ap_rst_n_Boundary_X4Y4_To_X6Y4_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper187_U0_fifo_w_out_V_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper187_U0_fifo_w_out_V_V_din_pass_1_q0 <= PE_wrapper187_U0_fifo_w_out_V_V_din_pass_1_out;
  end
  assign PE_wrapper187_U0_fifo_w_out_V_V_din_pass_1_in = PE_wrapper187_U0_fifo_w_out_V_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_3_2_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_3_2_V_V_full_n_pass_0_q0 <= fifo_w_PE_3_2_V_V_full_n_pass_0_out;
  end
  assign fifo_w_PE_3_2_V_V_full_n_pass_0_in = fifo_w_PE_3_2_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper187_U0_fifo_w_out_V_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper187_U0_fifo_w_out_V_V_write_pass_1_q0 <= PE_wrapper187_U0_fifo_w_out_V_V_write_pass_1_out;
  end
  assign PE_wrapper187_U0_fifo_w_out_V_V_write_pass_1_in = PE_wrapper187_U0_fifo_w_out_V_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [31:0] PE_wrapper163_U0_fifo_cout_drain_out_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper163_U0_fifo_cout_drain_out_V_din_pass_1_q0 <= PE_wrapper163_U0_fifo_cout_drain_out_V_din_pass_1_out;
  end
  assign PE_wrapper163_U0_fifo_cout_drain_out_V_din_pass_1_in = PE_wrapper163_U0_fifo_cout_drain_out_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_PE_1_1_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_PE_1_1_V_full_n_pass_0_q0 <= fifo_cout_drain_PE_1_1_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_PE_1_1_V_full_n_pass_0_in = fifo_cout_drain_PE_1_1_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper163_U0_fifo_cout_drain_out_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper163_U0_fifo_cout_drain_out_V_write_pass_1_q0 <= PE_wrapper163_U0_fifo_cout_drain_out_V_write_pass_1_out;
  end
  assign PE_wrapper163_U0_fifo_cout_drain_out_V_write_pass_1_in = PE_wrapper163_U0_fifo_cout_drain_out_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [31:0] PE_wrapper175_U0_fifo_cout_drain_out_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper175_U0_fifo_cout_drain_out_V_din_pass_1_q0 <= PE_wrapper175_U0_fifo_cout_drain_out_V_din_pass_1_out;
  end
  assign PE_wrapper175_U0_fifo_cout_drain_out_V_din_pass_1_in = PE_wrapper175_U0_fifo_cout_drain_out_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_PE_2_1_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_PE_2_1_V_full_n_pass_0_q0 <= fifo_cout_drain_PE_2_1_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_PE_2_1_V_full_n_pass_0_in = fifo_cout_drain_PE_2_1_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper175_U0_fifo_cout_drain_out_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper175_U0_fifo_cout_drain_out_V_write_pass_1_q0 <= PE_wrapper175_U0_fifo_cout_drain_out_V_write_pass_1_out;
  end
  assign PE_wrapper175_U0_fifo_cout_drain_out_V_write_pass_1_in = PE_wrapper175_U0_fifo_cout_drain_out_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper187_U0_fifo_cin_out_V_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper187_U0_fifo_cin_out_V_V_din_pass_1_q0 <= PE_wrapper187_U0_fifo_cin_out_V_V_din_pass_1_out;
  end
  assign PE_wrapper187_U0_fifo_cin_out_V_V_din_pass_1_in = PE_wrapper187_U0_fifo_cin_out_V_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_4_1_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_4_1_V_V_full_n_pass_0_q0 <= fifo_cin_PE_4_1_V_V_full_n_pass_0_out;
  end
  assign fifo_cin_PE_4_1_V_V_full_n_pass_0_in = fifo_cin_PE_4_1_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper187_U0_fifo_cin_out_V_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper187_U0_fifo_cin_out_V_V_write_pass_1_q0 <= PE_wrapper187_U0_fifo_cin_out_V_V_write_pass_1_out;
  end
  assign PE_wrapper187_U0_fifo_cin_out_V_V_write_pass_1_in = PE_wrapper187_U0_fifo_cin_out_V_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper186_U0_fifo_cin_out_V_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper186_U0_fifo_cin_out_V_V_din_pass_1_q0 <= PE_wrapper186_U0_fifo_cin_out_V_V_din_pass_1_out;
  end
  assign PE_wrapper186_U0_fifo_cin_out_V_V_din_pass_1_in = PE_wrapper186_U0_fifo_cin_out_V_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_4_0_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_4_0_V_V_full_n_pass_0_q0 <= fifo_cin_PE_4_0_V_V_full_n_pass_0_out;
  end
  assign fifo_cin_PE_4_0_V_V_full_n_pass_0_in = fifo_cin_PE_4_0_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper186_U0_fifo_cin_out_V_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper186_U0_fifo_cin_out_V_V_write_pass_1_q0 <= PE_wrapper186_U0_fifo_cin_out_V_V_write_pass_1_out;
  end
  assign PE_wrapper186_U0_fifo_cin_out_V_V_write_pass_1_in = PE_wrapper186_U0_fifo_cin_out_V_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [31:0] PE_wrapper187_U0_fifo_cout_drain_out_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper187_U0_fifo_cout_drain_out_V_din_pass_1_q0 <= PE_wrapper187_U0_fifo_cout_drain_out_V_din_pass_1_out;
  end
  assign PE_wrapper187_U0_fifo_cout_drain_out_V_din_pass_1_in = PE_wrapper187_U0_fifo_cout_drain_out_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_PE_3_1_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_PE_3_1_V_full_n_pass_0_q0 <= fifo_cout_drain_PE_3_1_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_PE_3_1_V_full_n_pass_0_in = fifo_cout_drain_PE_3_1_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper187_U0_fifo_cout_drain_out_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper187_U0_fifo_cout_drain_out_V_write_pass_1_q0 <= PE_wrapper187_U0_fifo_cout_drain_out_V_write_pass_1_out;
  end
  assign PE_wrapper187_U0_fifo_cout_drain_out_V_write_pass_1_in = PE_wrapper187_U0_fifo_cout_drain_out_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [255:0] w_IO_L2_in137_U0_fifo_w_out_V_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    w_IO_L2_in137_U0_fifo_w_out_V_V_din_pass_1_q0 <= w_IO_L2_in137_U0_fifo_w_out_V_V_din_pass_1_out;
  end
  assign w_IO_L2_in137_U0_fifo_w_out_V_V_din_pass_1_in = w_IO_L2_in137_U0_fifo_w_out_V_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_w_w_IO_L2_in_3_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_w_IO_L2_in_3_V_V_full_n_pass_0_q0 <= fifo_w_w_IO_L2_in_3_V_V_full_n_pass_0_out;
  end
  assign fifo_w_w_IO_L2_in_3_V_V_full_n_pass_0_in = fifo_w_w_IO_L2_in_3_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  w_IO_L2_in137_U0_fifo_w_out_V_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    w_IO_L2_in137_U0_fifo_w_out_V_V_write_pass_1_q0 <= w_IO_L2_in137_U0_fifo_w_out_V_V_write_pass_1_out;
  end
  assign w_IO_L2_in137_U0_fifo_w_out_V_V_write_pass_1_in = w_IO_L2_in137_U0_fifo_w_out_V_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [63:0] cout_drain_IO_L1_out_wrapper376_U0_fifo_cout_drain_out_V_V_din_pass_2_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper376_U0_fifo_cout_drain_out_V_V_din_pass_2_q0 <= cout_drain_IO_L1_out_wrapper376_U0_fifo_cout_drain_out_V_V_din_pass_2_out;
  end
  assign cout_drain_IO_L1_out_wrapper376_U0_fifo_cout_drain_out_V_V_din_pass_2_in = cout_drain_IO_L1_out_wrapper376_U0_fifo_cout_drain_out_V_V_din_pass_2_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_cout_drain_IO_L1_out_0_6_V_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_cout_drain_IO_L1_out_0_6_V_V_full_n_pass_1_q0 <= fifo_cout_drain_cout_drain_IO_L1_out_0_6_V_V_full_n_pass_1_out;
  end
  assign fifo_cout_drain_cout_drain_IO_L1_out_0_6_V_V_full_n_pass_1_in = fifo_cout_drain_cout_drain_IO_L1_out_0_6_V_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg  cout_drain_IO_L1_out_wrapper376_U0_fifo_cout_drain_out_V_V_write_pass_2_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper376_U0_fifo_cout_drain_out_V_V_write_pass_2_q0 <= cout_drain_IO_L1_out_wrapper376_U0_fifo_cout_drain_out_V_V_write_pass_2_out;
  end
  assign cout_drain_IO_L1_out_wrapper376_U0_fifo_cout_drain_out_V_V_write_pass_2_in = cout_drain_IO_L1_out_wrapper376_U0_fifo_cout_drain_out_V_V_write_pass_2_q0;
  (* dont_touch = "yes" *) reg [31:0] PE_wrapper151_U0_fifo_cout_drain_out_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper151_U0_fifo_cout_drain_out_V_din_pass_1_q0 <= PE_wrapper151_U0_fifo_cout_drain_out_V_din_pass_1_out;
  end
  assign PE_wrapper151_U0_fifo_cout_drain_out_V_din_pass_1_in = PE_wrapper151_U0_fifo_cout_drain_out_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_PE_0_1_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_PE_0_1_V_full_n_pass_0_q0 <= fifo_cout_drain_PE_0_1_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_PE_0_1_V_full_n_pass_0_in = fifo_cout_drain_PE_0_1_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper151_U0_fifo_cout_drain_out_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper151_U0_fifo_cout_drain_out_V_write_pass_1_q0 <= PE_wrapper151_U0_fifo_cout_drain_out_V_write_pass_1_out;
  end
  assign PE_wrapper151_U0_fifo_cout_drain_out_V_write_pass_1_in = PE_wrapper151_U0_fifo_cout_drain_out_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [63:0] cout_drain_IO_L1_out_wrapper392_U0_fifo_cout_drain_out_V_V_din_pass_2_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper392_U0_fifo_cout_drain_out_V_V_din_pass_2_q0 <= cout_drain_IO_L1_out_wrapper392_U0_fifo_cout_drain_out_V_V_din_pass_2_out;
  end
  assign cout_drain_IO_L1_out_wrapper392_U0_fifo_cout_drain_out_V_V_din_pass_2_in = cout_drain_IO_L1_out_wrapper392_U0_fifo_cout_drain_out_V_V_din_pass_2_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_cout_drain_IO_L1_out_1_6_V_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_cout_drain_IO_L1_out_1_6_V_V_full_n_pass_1_q0 <= fifo_cout_drain_cout_drain_IO_L1_out_1_6_V_V_full_n_pass_1_out;
  end
  assign fifo_cout_drain_cout_drain_IO_L1_out_1_6_V_V_full_n_pass_1_in = fifo_cout_drain_cout_drain_IO_L1_out_1_6_V_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg  cout_drain_IO_L1_out_wrapper392_U0_fifo_cout_drain_out_V_V_write_pass_2_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper392_U0_fifo_cout_drain_out_V_V_write_pass_2_q0 <= cout_drain_IO_L1_out_wrapper392_U0_fifo_cout_drain_out_V_V_write_pass_2_out;
  end
  assign cout_drain_IO_L1_out_wrapper392_U0_fifo_cout_drain_out_V_V_write_pass_2_in = cout_drain_IO_L1_out_wrapper392_U0_fifo_cout_drain_out_V_V_write_pass_2_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_cout_drain_IO_L2_out_4_V_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_cout_drain_IO_L2_out_4_V_V_full_n_pass_1_q0 <= fifo_cout_drain_cout_drain_IO_L2_out_4_V_V_full_n_pass_1_out;
  end
  assign fifo_cout_drain_cout_drain_IO_L2_out_4_V_V_full_n_pass_1_in = fifo_cout_drain_cout_drain_IO_L2_out_4_V_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_PE_4_2_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_PE_4_2_V_full_n_pass_0_q0 <= fifo_cout_drain_PE_4_2_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_PE_4_2_V_full_n_pass_0_in = fifo_cout_drain_PE_4_2_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper212_U0_fifo_cin_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper212_U0_fifo_cin_out_V_V_din_pass_0_q0 <= PE_wrapper212_U0_fifo_cin_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper212_U0_fifo_cin_out_V_V_din_pass_0_in = PE_wrapper212_U0_fifo_cin_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper212_U0_fifo_cin_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper212_U0_fifo_cin_out_V_V_write_pass_0_q0 <= PE_wrapper212_U0_fifo_cin_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper212_U0_fifo_cin_out_V_V_write_pass_0_in = PE_wrapper212_U0_fifo_cin_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_5_1_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_5_1_V_V_full_n_pass_0_q0 <= fifo_w_PE_5_1_V_V_full_n_pass_0_out;
  end
  assign fifo_w_PE_5_1_V_V_full_n_pass_0_in = fifo_w_PE_5_1_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_PE_3_2_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_PE_3_2_V_full_n_pass_0_q0 <= fifo_cout_drain_PE_3_2_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_PE_3_2_V_full_n_pass_0_in = fifo_cout_drain_PE_3_2_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_cout_drain_IO_L1_out_3_6_V_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_cout_drain_IO_L1_out_3_6_V_V_full_n_pass_1_q0 <= fifo_cout_drain_cout_drain_IO_L1_out_3_6_V_V_full_n_pass_1_out;
  end
  assign fifo_cout_drain_cout_drain_IO_L1_out_3_6_V_V_full_n_pass_1_in = fifo_cout_drain_cout_drain_IO_L1_out_3_6_V_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_5_3_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_5_3_V_V_full_n_pass_0_q0 <= fifo_cin_PE_5_3_V_V_full_n_pass_0_out;
  end
  assign fifo_cin_PE_5_3_V_V_full_n_pass_0_in = fifo_cin_PE_5_3_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_cout_drain_IO_L1_out_1_0_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_cout_drain_IO_L1_out_1_0_V_V_full_n_pass_0_q0 <= fifo_cout_drain_cout_drain_IO_L1_out_1_0_V_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_cout_drain_IO_L1_out_1_0_V_V_full_n_pass_0_in = fifo_cout_drain_cout_drain_IO_L1_out_1_0_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_5_1_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_5_1_V_V_full_n_pass_0_q0 <= fifo_cin_PE_5_1_V_V_full_n_pass_0_out;
  end
  assign fifo_cin_PE_5_1_V_V_full_n_pass_0_in = fifo_cin_PE_5_1_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper211_U0_fifo_cin_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper211_U0_fifo_cin_out_V_V_din_pass_0_q0 <= PE_wrapper211_U0_fifo_cin_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper211_U0_fifo_cin_out_V_V_din_pass_0_in = PE_wrapper211_U0_fifo_cin_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper211_U0_fifo_cin_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper211_U0_fifo_cin_out_V_V_write_pass_0_q0 <= PE_wrapper211_U0_fifo_cin_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper211_U0_fifo_cin_out_V_V_write_pass_0_in = PE_wrapper211_U0_fifo_cin_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_PE_1_3_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_PE_1_3_V_full_n_pass_1_q0 <= fifo_cout_drain_PE_1_3_V_full_n_pass_1_out;
  end
  assign fifo_cout_drain_PE_1_3_V_full_n_pass_1_in = fifo_cout_drain_PE_1_3_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg [31:0] PE_wrapper211_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper211_U0_fifo_cout_drain_out_V_din_pass_0_q0 <= PE_wrapper211_U0_fifo_cout_drain_out_V_din_pass_0_out;
  end
  assign PE_wrapper211_U0_fifo_cout_drain_out_V_din_pass_0_in = PE_wrapper211_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper211_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper211_U0_fifo_cout_drain_out_V_write_pass_0_q0 <= PE_wrapper211_U0_fifo_cout_drain_out_V_write_pass_0_out;
  end
  assign PE_wrapper211_U0_fifo_cout_drain_out_V_write_pass_0_in = PE_wrapper211_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_PE_0_3_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_PE_0_3_V_full_n_pass_1_q0 <= fifo_cout_drain_PE_0_3_V_full_n_pass_1_out;
  end
  assign fifo_cout_drain_PE_0_3_V_full_n_pass_1_in = fifo_cout_drain_PE_0_3_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_PE_4_3_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_PE_4_3_V_full_n_pass_0_q0 <= fifo_cout_drain_PE_4_3_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_PE_4_3_V_full_n_pass_0_in = fifo_cout_drain_PE_4_3_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_cout_drain_IO_L1_out_0_0_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_cout_drain_IO_L1_out_0_0_V_V_full_n_pass_0_q0 <= fifo_cout_drain_cout_drain_IO_L1_out_0_0_V_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_cout_drain_IO_L1_out_0_0_V_V_full_n_pass_0_in = fifo_cout_drain_cout_drain_IO_L1_out_0_0_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper213_U0_fifo_cin_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper213_U0_fifo_cin_out_V_V_din_pass_0_q0 <= PE_wrapper213_U0_fifo_cin_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper213_U0_fifo_cin_out_V_V_din_pass_0_in = PE_wrapper213_U0_fifo_cin_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper213_U0_fifo_cin_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper213_U0_fifo_cin_out_V_V_write_pass_0_q0 <= PE_wrapper213_U0_fifo_cin_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper213_U0_fifo_cin_out_V_V_write_pass_0_in = PE_wrapper213_U0_fifo_cin_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_PE_2_3_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_PE_2_3_V_full_n_pass_1_q0 <= fifo_cout_drain_PE_2_3_V_full_n_pass_1_out;
  end
  assign fifo_cout_drain_PE_2_3_V_full_n_pass_1_in = fifo_cout_drain_PE_2_3_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_PE_1_2_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_PE_1_2_V_full_n_pass_1_q0 <= fifo_cout_drain_PE_1_2_V_full_n_pass_1_out;
  end
  assign fifo_cout_drain_PE_1_2_V_full_n_pass_1_in = fifo_cout_drain_PE_1_2_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_PE_3_3_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_PE_3_3_V_full_n_pass_1_q0 <= fifo_cout_drain_PE_3_3_V_full_n_pass_1_out;
  end
  assign fifo_cout_drain_PE_3_3_V_full_n_pass_1_in = fifo_cout_drain_PE_3_3_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_cin_IO_L2_in_1_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_cin_IO_L2_in_1_V_V_full_n_pass_0_q0 <= fifo_cin_cin_IO_L2_in_1_V_V_full_n_pass_0_out;
  end
  assign fifo_cin_cin_IO_L2_in_1_V_V_full_n_pass_0_in = fifo_cin_cin_IO_L2_in_1_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_PE_0_2_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_PE_0_2_V_full_n_pass_1_q0 <= fifo_cout_drain_PE_0_2_V_full_n_pass_1_out;
  end
  assign fifo_cout_drain_PE_0_2_V_full_n_pass_1_in = fifo_cout_drain_PE_0_2_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg [255:0] cin_IO_L2_in125_U0_fifo_cin_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    cin_IO_L2_in125_U0_fifo_cin_out_V_V_din_pass_0_q0 <= cin_IO_L2_in125_U0_fifo_cin_out_V_V_din_pass_0_out;
  end
  assign cin_IO_L2_in125_U0_fifo_cin_out_V_V_din_pass_0_in = cin_IO_L2_in125_U0_fifo_cin_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  cin_IO_L2_in125_U0_fifo_cin_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    cin_IO_L2_in125_U0_fifo_cin_out_V_V_write_pass_0_q0 <= cin_IO_L2_in125_U0_fifo_cin_out_V_V_write_pass_0_out;
  end
  assign cin_IO_L2_in125_U0_fifo_cin_out_V_V_write_pass_0_in = cin_IO_L2_in125_U0_fifo_cin_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_5_2_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_5_2_V_V_full_n_pass_0_q0 <= fifo_cin_PE_5_2_V_V_full_n_pass_0_out;
  end
  assign fifo_cin_PE_5_2_V_V_full_n_pass_0_in = fifo_cin_PE_5_2_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] cin_IO_L2_in125_U0_fifo_cin_local_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    cin_IO_L2_in125_U0_fifo_cin_local_out_V_V_din_pass_0_q0 <= cin_IO_L2_in125_U0_fifo_cin_local_out_V_V_din_pass_0_out;
  end
  assign cin_IO_L2_in125_U0_fifo_cin_local_out_V_V_din_pass_0_in = cin_IO_L2_in125_U0_fifo_cin_local_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  cin_IO_L2_in125_U0_fifo_cin_local_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    cin_IO_L2_in125_U0_fifo_cin_local_out_V_V_write_pass_0_q0 <= cin_IO_L2_in125_U0_fifo_cin_local_out_V_V_write_pass_0_out;
  end
  assign cin_IO_L2_in125_U0_fifo_cin_local_out_V_V_write_pass_0_in = cin_IO_L2_in125_U0_fifo_cin_local_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_cout_drain_IO_L1_out_2_6_V_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_cout_drain_IO_L1_out_2_6_V_V_full_n_pass_1_q0 <= fifo_cout_drain_cout_drain_IO_L1_out_2_6_V_V_full_n_pass_1_out;
  end
  assign fifo_cout_drain_cout_drain_IO_L1_out_2_6_V_V_full_n_pass_1_in = fifo_cout_drain_cout_drain_IO_L1_out_2_6_V_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper213_U0_fifo_w_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper213_U0_fifo_w_out_V_V_din_pass_0_q0 <= PE_wrapper213_U0_fifo_w_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper213_U0_fifo_w_out_V_V_din_pass_0_in = PE_wrapper213_U0_fifo_w_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper213_U0_fifo_w_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper213_U0_fifo_w_out_V_V_write_pass_0_q0 <= PE_wrapper213_U0_fifo_w_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper213_U0_fifo_w_out_V_V_write_pass_0_in = PE_wrapper213_U0_fifo_w_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [63:0] cout_drain_IO_L2_out568_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L2_out568_U0_fifo_cout_drain_out_V_V_din_pass_0_q0 <= cout_drain_IO_L2_out568_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  end
  assign cout_drain_IO_L2_out568_U0_fifo_cout_drain_out_V_V_din_pass_0_in = cout_drain_IO_L2_out568_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  cout_drain_IO_L2_out568_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L2_out568_U0_fifo_cout_drain_out_V_V_write_pass_0_q0 <= cout_drain_IO_L2_out568_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  end
  assign cout_drain_IO_L2_out568_U0_fifo_cout_drain_out_V_V_write_pass_0_in = cout_drain_IO_L2_out568_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_PE_2_2_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_PE_2_2_V_full_n_pass_1_q0 <= fifo_cout_drain_PE_2_2_V_full_n_pass_1_out;
  end
  assign fifo_cout_drain_PE_2_2_V_full_n_pass_1_in = fifo_cout_drain_PE_2_2_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg  ap_done_Boundary_X6Y0_To_X6Y2_q0;
  always @ (posedge ap_clk) begin
    ap_done_Boundary_X6Y0_To_X6Y2_q0 <= ap_done_Boundary_X6Y0_To_X6Y2_out;
  end
  assign ap_done_Boundary_X6Y0_To_X6Y2_in = ap_done_Boundary_X6Y0_To_X6Y2_q0;
  (* dont_touch = "yes" *) reg  ap_start_Boundary_X6Y2_To_X8Y2_q0;
  always @ (posedge ap_clk) begin
    ap_start_Boundary_X6Y2_To_X8Y2_q0 <= ap_start_Boundary_X6Y2_To_X8Y2_out;
  end
  assign ap_start_Boundary_X6Y2_To_X8Y2_in = ap_start_Boundary_X6Y2_To_X8Y2_q0;
  (* dont_touch = "yes" *) reg  ap_rst_n_Boundary_X6Y2_To_X8Y2_q0;
  always @ (posedge ap_clk) begin
    ap_rst_n_Boundary_X6Y2_To_X8Y2_q0 <= ap_rst_n_Boundary_X6Y2_To_X8Y2_out;
  end
  assign ap_rst_n_Boundary_X6Y2_To_X8Y2_in = ap_rst_n_Boundary_X6Y2_To_X8Y2_q0;
  (* dont_touch = "yes" *) reg [63:0] cout_drain_IO_L2_out564_U0_fifo_cout_drain_out_V_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L2_out564_U0_fifo_cout_drain_out_V_V_din_pass_1_q0 <= cout_drain_IO_L2_out564_U0_fifo_cout_drain_out_V_V_din_pass_1_out;
  end
  assign cout_drain_IO_L2_out564_U0_fifo_cout_drain_out_V_V_din_pass_1_in = cout_drain_IO_L2_out564_U0_fifo_cout_drain_out_V_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_cout_drain_IO_L2_out_4_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_cout_drain_IO_L2_out_4_V_V_full_n_pass_0_q0 <= fifo_cout_drain_cout_drain_IO_L2_out_4_V_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_cout_drain_IO_L2_out_4_V_V_full_n_pass_0_in = fifo_cout_drain_cout_drain_IO_L2_out_4_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  cout_drain_IO_L2_out564_U0_fifo_cout_drain_out_V_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L2_out564_U0_fifo_cout_drain_out_V_V_write_pass_1_q0 <= cout_drain_IO_L2_out564_U0_fifo_cout_drain_out_V_V_write_pass_1_out;
  end
  assign cout_drain_IO_L2_out564_U0_fifo_cout_drain_out_V_V_write_pass_1_in = cout_drain_IO_L2_out564_U0_fifo_cout_drain_out_V_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [31:0] PE_wrapper165_U0_fifo_cout_drain_out_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper165_U0_fifo_cout_drain_out_V_din_pass_1_q0 <= PE_wrapper165_U0_fifo_cout_drain_out_V_din_pass_1_out;
  end
  assign PE_wrapper165_U0_fifo_cout_drain_out_V_din_pass_1_in = PE_wrapper165_U0_fifo_cout_drain_out_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_PE_1_3_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_PE_1_3_V_full_n_pass_0_q0 <= fifo_cout_drain_PE_1_3_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_PE_1_3_V_full_n_pass_0_in = fifo_cout_drain_PE_1_3_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper165_U0_fifo_cout_drain_out_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper165_U0_fifo_cout_drain_out_V_write_pass_1_q0 <= PE_wrapper165_U0_fifo_cout_drain_out_V_write_pass_1_out;
  end
  assign PE_wrapper165_U0_fifo_cout_drain_out_V_write_pass_1_in = PE_wrapper165_U0_fifo_cout_drain_out_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [31:0] PE_wrapper153_U0_fifo_cout_drain_out_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper153_U0_fifo_cout_drain_out_V_din_pass_1_q0 <= PE_wrapper153_U0_fifo_cout_drain_out_V_din_pass_1_out;
  end
  assign PE_wrapper153_U0_fifo_cout_drain_out_V_din_pass_1_in = PE_wrapper153_U0_fifo_cout_drain_out_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_PE_0_3_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_PE_0_3_V_full_n_pass_0_q0 <= fifo_cout_drain_PE_0_3_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_PE_0_3_V_full_n_pass_0_in = fifo_cout_drain_PE_0_3_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper153_U0_fifo_cout_drain_out_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper153_U0_fifo_cout_drain_out_V_write_pass_1_q0 <= PE_wrapper153_U0_fifo_cout_drain_out_V_write_pass_1_out;
  end
  assign PE_wrapper153_U0_fifo_cout_drain_out_V_write_pass_1_in = PE_wrapper153_U0_fifo_cout_drain_out_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [31:0] PE_wrapper177_U0_fifo_cout_drain_out_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper177_U0_fifo_cout_drain_out_V_din_pass_1_q0 <= PE_wrapper177_U0_fifo_cout_drain_out_V_din_pass_1_out;
  end
  assign PE_wrapper177_U0_fifo_cout_drain_out_V_din_pass_1_in = PE_wrapper177_U0_fifo_cout_drain_out_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_PE_2_3_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_PE_2_3_V_full_n_pass_0_q0 <= fifo_cout_drain_PE_2_3_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_PE_2_3_V_full_n_pass_0_in = fifo_cout_drain_PE_2_3_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper177_U0_fifo_cout_drain_out_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper177_U0_fifo_cout_drain_out_V_write_pass_1_q0 <= PE_wrapper177_U0_fifo_cout_drain_out_V_write_pass_1_out;
  end
  assign PE_wrapper177_U0_fifo_cout_drain_out_V_write_pass_1_in = PE_wrapper177_U0_fifo_cout_drain_out_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [31:0] PE_wrapper164_U0_fifo_cout_drain_out_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper164_U0_fifo_cout_drain_out_V_din_pass_1_q0 <= PE_wrapper164_U0_fifo_cout_drain_out_V_din_pass_1_out;
  end
  assign PE_wrapper164_U0_fifo_cout_drain_out_V_din_pass_1_in = PE_wrapper164_U0_fifo_cout_drain_out_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_PE_1_2_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_PE_1_2_V_full_n_pass_0_q0 <= fifo_cout_drain_PE_1_2_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_PE_1_2_V_full_n_pass_0_in = fifo_cout_drain_PE_1_2_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper164_U0_fifo_cout_drain_out_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper164_U0_fifo_cout_drain_out_V_write_pass_1_q0 <= PE_wrapper164_U0_fifo_cout_drain_out_V_write_pass_1_out;
  end
  assign PE_wrapper164_U0_fifo_cout_drain_out_V_write_pass_1_in = PE_wrapper164_U0_fifo_cout_drain_out_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [31:0] PE_wrapper189_U0_fifo_cout_drain_out_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper189_U0_fifo_cout_drain_out_V_din_pass_1_q0 <= PE_wrapper189_U0_fifo_cout_drain_out_V_din_pass_1_out;
  end
  assign PE_wrapper189_U0_fifo_cout_drain_out_V_din_pass_1_in = PE_wrapper189_U0_fifo_cout_drain_out_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_PE_3_3_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_PE_3_3_V_full_n_pass_0_q0 <= fifo_cout_drain_PE_3_3_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_PE_3_3_V_full_n_pass_0_in = fifo_cout_drain_PE_3_3_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper189_U0_fifo_cout_drain_out_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper189_U0_fifo_cout_drain_out_V_write_pass_1_q0 <= PE_wrapper189_U0_fifo_cout_drain_out_V_write_pass_1_out;
  end
  assign PE_wrapper189_U0_fifo_cout_drain_out_V_write_pass_1_in = PE_wrapper189_U0_fifo_cout_drain_out_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [31:0] PE_wrapper152_U0_fifo_cout_drain_out_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper152_U0_fifo_cout_drain_out_V_din_pass_1_q0 <= PE_wrapper152_U0_fifo_cout_drain_out_V_din_pass_1_out;
  end
  assign PE_wrapper152_U0_fifo_cout_drain_out_V_din_pass_1_in = PE_wrapper152_U0_fifo_cout_drain_out_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_PE_0_2_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_PE_0_2_V_full_n_pass_0_q0 <= fifo_cout_drain_PE_0_2_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_PE_0_2_V_full_n_pass_0_in = fifo_cout_drain_PE_0_2_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper152_U0_fifo_cout_drain_out_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper152_U0_fifo_cout_drain_out_V_write_pass_1_q0 <= PE_wrapper152_U0_fifo_cout_drain_out_V_write_pass_1_out;
  end
  assign PE_wrapper152_U0_fifo_cout_drain_out_V_write_pass_1_in = PE_wrapper152_U0_fifo_cout_drain_out_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [31:0] PE_wrapper176_U0_fifo_cout_drain_out_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper176_U0_fifo_cout_drain_out_V_din_pass_1_q0 <= PE_wrapper176_U0_fifo_cout_drain_out_V_din_pass_1_out;
  end
  assign PE_wrapper176_U0_fifo_cout_drain_out_V_din_pass_1_in = PE_wrapper176_U0_fifo_cout_drain_out_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_PE_2_2_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_PE_2_2_V_full_n_pass_0_q0 <= fifo_cout_drain_PE_2_2_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_PE_2_2_V_full_n_pass_0_in = fifo_cout_drain_PE_2_2_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper176_U0_fifo_cout_drain_out_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper176_U0_fifo_cout_drain_out_V_write_pass_1_q0 <= PE_wrapper176_U0_fifo_cout_drain_out_V_write_pass_1_out;
  end
  assign PE_wrapper176_U0_fifo_cout_drain_out_V_write_pass_1_in = PE_wrapper176_U0_fifo_cout_drain_out_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper165_U0_fifo_w_out_V_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper165_U0_fifo_w_out_V_V_din_pass_1_q0 <= PE_wrapper165_U0_fifo_w_out_V_V_din_pass_1_out;
  end
  assign PE_wrapper165_U0_fifo_w_out_V_V_din_pass_1_in = PE_wrapper165_U0_fifo_w_out_V_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_1_4_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_1_4_V_V_full_n_pass_0_q0 <= fifo_w_PE_1_4_V_V_full_n_pass_0_out;
  end
  assign fifo_w_PE_1_4_V_V_full_n_pass_0_in = fifo_w_PE_1_4_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper165_U0_fifo_w_out_V_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper165_U0_fifo_w_out_V_V_write_pass_1_q0 <= PE_wrapper165_U0_fifo_w_out_V_V_write_pass_1_out;
  end
  assign PE_wrapper165_U0_fifo_w_out_V_V_write_pass_1_in = PE_wrapper165_U0_fifo_w_out_V_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [255:0] cin_IO_L2_in127_U0_fifo_cin_out_V_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    cin_IO_L2_in127_U0_fifo_cin_out_V_V_din_pass_1_q0 <= cin_IO_L2_in127_U0_fifo_cin_out_V_V_din_pass_1_out;
  end
  assign cin_IO_L2_in127_U0_fifo_cin_out_V_V_din_pass_1_in = cin_IO_L2_in127_U0_fifo_cin_out_V_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_cin_IO_L2_in_4_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_cin_IO_L2_in_4_V_V_full_n_pass_0_q0 <= fifo_cin_cin_IO_L2_in_4_V_V_full_n_pass_0_out;
  end
  assign fifo_cin_cin_IO_L2_in_4_V_V_full_n_pass_0_in = fifo_cin_cin_IO_L2_in_4_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  cin_IO_L2_in127_U0_fifo_cin_out_V_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    cin_IO_L2_in127_U0_fifo_cin_out_V_V_write_pass_1_q0 <= cin_IO_L2_in127_U0_fifo_cin_out_V_V_write_pass_1_out;
  end
  assign cin_IO_L2_in127_U0_fifo_cin_out_V_V_write_pass_1_in = cin_IO_L2_in127_U0_fifo_cin_out_V_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper177_U0_fifo_w_out_V_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper177_U0_fifo_w_out_V_V_din_pass_1_q0 <= PE_wrapper177_U0_fifo_w_out_V_V_din_pass_1_out;
  end
  assign PE_wrapper177_U0_fifo_w_out_V_V_din_pass_1_in = PE_wrapper177_U0_fifo_w_out_V_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_2_4_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_2_4_V_V_full_n_pass_0_q0 <= fifo_w_PE_2_4_V_V_full_n_pass_0_out;
  end
  assign fifo_w_PE_2_4_V_V_full_n_pass_0_in = fifo_w_PE_2_4_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper177_U0_fifo_w_out_V_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper177_U0_fifo_w_out_V_V_write_pass_1_q0 <= PE_wrapper177_U0_fifo_w_out_V_V_write_pass_1_out;
  end
  assign PE_wrapper177_U0_fifo_w_out_V_V_write_pass_1_in = PE_wrapper177_U0_fifo_w_out_V_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper153_U0_fifo_w_out_V_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper153_U0_fifo_w_out_V_V_din_pass_1_q0 <= PE_wrapper153_U0_fifo_w_out_V_V_din_pass_1_out;
  end
  assign PE_wrapper153_U0_fifo_w_out_V_V_din_pass_1_in = PE_wrapper153_U0_fifo_w_out_V_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_0_4_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_0_4_V_V_full_n_pass_0_q0 <= fifo_w_PE_0_4_V_V_full_n_pass_0_out;
  end
  assign fifo_w_PE_0_4_V_V_full_n_pass_0_in = fifo_w_PE_0_4_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper153_U0_fifo_w_out_V_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper153_U0_fifo_w_out_V_V_write_pass_1_q0 <= PE_wrapper153_U0_fifo_w_out_V_V_write_pass_1_out;
  end
  assign PE_wrapper153_U0_fifo_w_out_V_V_write_pass_1_in = PE_wrapper153_U0_fifo_w_out_V_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper189_U0_fifo_w_out_V_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper189_U0_fifo_w_out_V_V_din_pass_1_q0 <= PE_wrapper189_U0_fifo_w_out_V_V_din_pass_1_out;
  end
  assign PE_wrapper189_U0_fifo_w_out_V_V_din_pass_1_in = PE_wrapper189_U0_fifo_w_out_V_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_3_4_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_3_4_V_V_full_n_pass_0_q0 <= fifo_w_PE_3_4_V_V_full_n_pass_0_out;
  end
  assign fifo_w_PE_3_4_V_V_full_n_pass_0_in = fifo_w_PE_3_4_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper189_U0_fifo_w_out_V_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper189_U0_fifo_w_out_V_V_write_pass_1_q0 <= PE_wrapper189_U0_fifo_w_out_V_V_write_pass_1_out;
  end
  assign PE_wrapper189_U0_fifo_w_out_V_V_write_pass_1_in = PE_wrapper189_U0_fifo_w_out_V_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [63:0] cout_drain_IO_L2_out568_U0_fifo_cout_drain_out_V_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L2_out568_U0_fifo_cout_drain_out_V_V_din_pass_1_q0 <= cout_drain_IO_L2_out568_U0_fifo_cout_drain_out_V_V_din_pass_1_out;
  end
  assign cout_drain_IO_L2_out568_U0_fifo_cout_drain_out_V_V_din_pass_1_in = cout_drain_IO_L2_out568_U0_fifo_cout_drain_out_V_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_cout_drain_IO_L2_out_0_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_cout_drain_IO_L2_out_0_V_V_full_n_pass_0_q0 <= fifo_cout_drain_cout_drain_IO_L2_out_0_V_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_cout_drain_IO_L2_out_0_V_V_full_n_pass_0_in = fifo_cout_drain_cout_drain_IO_L2_out_0_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  cout_drain_IO_L2_out568_U0_fifo_cout_drain_out_V_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L2_out568_U0_fifo_cout_drain_out_V_V_write_pass_1_q0 <= cout_drain_IO_L2_out568_U0_fifo_cout_drain_out_V_V_write_pass_1_out;
  end
  assign cout_drain_IO_L2_out568_U0_fifo_cout_drain_out_V_V_write_pass_1_in = cout_drain_IO_L2_out568_U0_fifo_cout_drain_out_V_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [255:0] w_IO_L2_in140_U0_fifo_w_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    w_IO_L2_in140_U0_fifo_w_out_V_V_din_pass_0_q0 <= w_IO_L2_in140_U0_fifo_w_out_V_V_din_pass_0_out;
  end
  assign w_IO_L2_in140_U0_fifo_w_out_V_V_din_pass_0_in = w_IO_L2_in140_U0_fifo_w_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  w_IO_L2_in140_U0_fifo_w_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    w_IO_L2_in140_U0_fifo_w_out_V_V_write_pass_0_q0 <= w_IO_L2_in140_U0_fifo_w_out_V_V_write_pass_0_out;
  end
  assign w_IO_L2_in140_U0_fifo_w_out_V_V_write_pass_0_in = w_IO_L2_in140_U0_fifo_w_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_3_2_V_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_3_2_V_V_full_n_pass_1_q0 <= fifo_w_PE_3_2_V_V_full_n_pass_1_out;
  end
  assign fifo_w_PE_3_2_V_V_full_n_pass_1_in = fifo_w_PE_3_2_V_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper188_U0_fifo_w_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper188_U0_fifo_w_out_V_V_din_pass_0_q0 <= PE_wrapper188_U0_fifo_w_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper188_U0_fifo_w_out_V_V_din_pass_0_in = PE_wrapper188_U0_fifo_w_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper188_U0_fifo_w_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper188_U0_fifo_w_out_V_V_write_pass_0_q0 <= PE_wrapper188_U0_fifo_w_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper188_U0_fifo_w_out_V_V_write_pass_0_in = PE_wrapper188_U0_fifo_w_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [31:0] PE_wrapper200_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper200_U0_fifo_cout_drain_out_V_din_pass_0_q0 <= PE_wrapper200_U0_fifo_cout_drain_out_V_din_pass_0_out;
  end
  assign PE_wrapper200_U0_fifo_cout_drain_out_V_din_pass_0_in = PE_wrapper200_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper200_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper200_U0_fifo_cout_drain_out_V_write_pass_0_q0 <= PE_wrapper200_U0_fifo_cout_drain_out_V_write_pass_0_out;
  end
  assign PE_wrapper200_U0_fifo_cout_drain_out_V_write_pass_0_in = PE_wrapper200_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [31:0] PE_wrapper188_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper188_U0_fifo_cout_drain_out_V_din_pass_0_q0 <= PE_wrapper188_U0_fifo_cout_drain_out_V_din_pass_0_out;
  end
  assign PE_wrapper188_U0_fifo_cout_drain_out_V_din_pass_0_in = PE_wrapper188_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper188_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper188_U0_fifo_cout_drain_out_V_write_pass_0_q0 <= PE_wrapper188_U0_fifo_cout_drain_out_V_write_pass_0_out;
  end
  assign PE_wrapper188_U0_fifo_cout_drain_out_V_write_pass_0_in = PE_wrapper188_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper210_U0_fifo_w_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper210_U0_fifo_w_out_V_V_din_pass_0_q0 <= PE_wrapper210_U0_fifo_w_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper210_U0_fifo_w_out_V_V_din_pass_0_in = PE_wrapper210_U0_fifo_w_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper210_U0_fifo_w_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper210_U0_fifo_w_out_V_V_write_pass_0_q0 <= PE_wrapper210_U0_fifo_w_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper210_U0_fifo_w_out_V_V_write_pass_0_in = PE_wrapper210_U0_fifo_w_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper201_U0_fifo_cin_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper201_U0_fifo_cin_out_V_V_din_pass_0_q0 <= PE_wrapper201_U0_fifo_cin_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper201_U0_fifo_cin_out_V_V_din_pass_0_in = PE_wrapper201_U0_fifo_cin_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper201_U0_fifo_cin_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper201_U0_fifo_cin_out_V_V_write_pass_0_q0 <= PE_wrapper201_U0_fifo_cin_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper201_U0_fifo_cin_out_V_V_write_pass_0_in = PE_wrapper201_U0_fifo_cin_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [63:0] cout_drain_IO_L1_out_wrapper398_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper398_U0_fifo_cout_drain_out_V_V_din_pass_0_q0 <= cout_drain_IO_L1_out_wrapper398_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper398_U0_fifo_cout_drain_out_V_V_din_pass_0_in = cout_drain_IO_L1_out_wrapper398_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  cout_drain_IO_L1_out_wrapper398_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper398_U0_fifo_cout_drain_out_V_V_write_pass_0_q0 <= cout_drain_IO_L1_out_wrapper398_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper398_U0_fifo_cout_drain_out_V_V_write_pass_0_in = cout_drain_IO_L1_out_wrapper398_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper199_U0_fifo_cin_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper199_U0_fifo_cin_out_V_V_din_pass_0_q0 <= PE_wrapper199_U0_fifo_cin_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper199_U0_fifo_cin_out_V_V_din_pass_0_in = PE_wrapper199_U0_fifo_cin_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper199_U0_fifo_cin_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper199_U0_fifo_cin_out_V_V_write_pass_0_q0 <= PE_wrapper199_U0_fifo_cin_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper199_U0_fifo_cin_out_V_V_write_pass_0_in = PE_wrapper199_U0_fifo_cin_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_PE_1_1_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_PE_1_1_V_full_n_pass_1_q0 <= fifo_cout_drain_PE_1_1_V_full_n_pass_1_out;
  end
  assign fifo_cout_drain_PE_1_1_V_full_n_pass_1_in = fifo_cout_drain_PE_1_1_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_PE_5_1_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_PE_5_1_V_full_n_pass_0_q0 <= fifo_cout_drain_PE_5_1_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_PE_5_1_V_full_n_pass_0_in = fifo_cout_drain_PE_5_1_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg [63:0] cout_drain_IO_L1_out_wrapper378_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper378_U0_fifo_cout_drain_out_V_V_din_pass_0_q0 <= cout_drain_IO_L1_out_wrapper378_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper378_U0_fifo_cout_drain_out_V_V_din_pass_0_in = cout_drain_IO_L1_out_wrapper378_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  cout_drain_IO_L1_out_wrapper378_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper378_U0_fifo_cout_drain_out_V_V_write_pass_0_q0 <= cout_drain_IO_L1_out_wrapper378_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper378_U0_fifo_cout_drain_out_V_V_write_pass_0_in = cout_drain_IO_L1_out_wrapper378_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_PE_2_1_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_PE_2_1_V_full_n_pass_1_q0 <= fifo_cout_drain_PE_2_1_V_full_n_pass_1_out;
  end
  assign fifo_cout_drain_PE_2_1_V_full_n_pass_1_in = fifo_cout_drain_PE_2_1_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg [31:0] PE_wrapper201_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper201_U0_fifo_cout_drain_out_V_din_pass_0_q0 <= PE_wrapper201_U0_fifo_cout_drain_out_V_din_pass_0_out;
  end
  assign PE_wrapper201_U0_fifo_cout_drain_out_V_din_pass_0_in = PE_wrapper201_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper201_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper201_U0_fifo_cout_drain_out_V_write_pass_0_q0 <= PE_wrapper201_U0_fifo_cout_drain_out_V_write_pass_0_out;
  end
  assign PE_wrapper201_U0_fifo_cout_drain_out_V_write_pass_0_in = PE_wrapper201_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_4_1_V_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_4_1_V_V_full_n_pass_1_q0 <= fifo_cin_PE_4_1_V_V_full_n_pass_1_out;
  end
  assign fifo_cin_PE_4_1_V_V_full_n_pass_1_in = fifo_cin_PE_4_1_V_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_4_0_V_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_4_0_V_V_full_n_pass_1_q0 <= fifo_cin_PE_4_0_V_V_full_n_pass_1_out;
  end
  assign fifo_cin_PE_4_0_V_V_full_n_pass_1_in = fifo_cin_PE_4_0_V_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper201_U0_fifo_w_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper201_U0_fifo_w_out_V_V_din_pass_0_q0 <= PE_wrapper201_U0_fifo_w_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper201_U0_fifo_w_out_V_V_din_pass_0_in = PE_wrapper201_U0_fifo_w_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper201_U0_fifo_w_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper201_U0_fifo_w_out_V_V_write_pass_0_q0 <= PE_wrapper201_U0_fifo_w_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper201_U0_fifo_w_out_V_V_write_pass_0_in = PE_wrapper201_U0_fifo_w_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_PE_3_1_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_PE_3_1_V_full_n_pass_1_q0 <= fifo_cout_drain_PE_3_1_V_full_n_pass_1_out;
  end
  assign fifo_cout_drain_PE_3_1_V_full_n_pass_1_in = fifo_cout_drain_PE_3_1_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_w_w_IO_L2_in_3_V_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_w_w_IO_L2_in_3_V_V_full_n_pass_1_q0 <= fifo_w_w_IO_L2_in_3_V_V_full_n_pass_1_out;
  end
  assign fifo_w_w_IO_L2_in_3_V_V_full_n_pass_1_in = fifo_w_w_IO_L2_in_3_V_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_cout_drain_IO_L1_out_0_6_V_V_full_n_pass_2_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_cout_drain_IO_L1_out_0_6_V_V_full_n_pass_2_q0 <= fifo_cout_drain_cout_drain_IO_L1_out_0_6_V_V_full_n_pass_2_out;
  end
  assign fifo_cout_drain_cout_drain_IO_L1_out_0_6_V_V_full_n_pass_2_in = fifo_cout_drain_cout_drain_IO_L1_out_0_6_V_V_full_n_pass_2_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_PE_0_1_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_PE_0_1_V_full_n_pass_1_q0 <= fifo_cout_drain_PE_0_1_V_full_n_pass_1_out;
  end
  assign fifo_cout_drain_PE_0_1_V_full_n_pass_1_in = fifo_cout_drain_PE_0_1_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg [255:0] w_IO_L2_in138_U0_fifo_w_local_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    w_IO_L2_in138_U0_fifo_w_local_out_V_V_din_pass_0_q0 <= w_IO_L2_in138_U0_fifo_w_local_out_V_V_din_pass_0_out;
  end
  assign w_IO_L2_in138_U0_fifo_w_local_out_V_V_din_pass_0_in = w_IO_L2_in138_U0_fifo_w_local_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  w_IO_L2_in138_U0_fifo_w_local_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    w_IO_L2_in138_U0_fifo_w_local_out_V_V_write_pass_0_q0 <= w_IO_L2_in138_U0_fifo_w_local_out_V_V_write_pass_0_out;
  end
  assign w_IO_L2_in138_U0_fifo_w_local_out_V_V_write_pass_0_in = w_IO_L2_in138_U0_fifo_w_local_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper200_U0_fifo_cin_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper200_U0_fifo_cin_out_V_V_din_pass_0_q0 <= PE_wrapper200_U0_fifo_cin_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper200_U0_fifo_cin_out_V_V_din_pass_0_in = PE_wrapper200_U0_fifo_cin_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper200_U0_fifo_cin_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper200_U0_fifo_cin_out_V_V_write_pass_0_q0 <= PE_wrapper200_U0_fifo_cin_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper200_U0_fifo_cin_out_V_V_write_pass_0_in = PE_wrapper200_U0_fifo_cin_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_4_3_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_4_3_V_V_full_n_pass_0_q0 <= fifo_cin_PE_4_3_V_V_full_n_pass_0_out;
  end
  assign fifo_cin_PE_4_3_V_V_full_n_pass_0_in = fifo_cin_PE_4_3_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_3_2_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_3_2_V_V_full_n_pass_0_q0 <= fifo_cin_PE_3_2_V_V_full_n_pass_0_out;
  end
  assign fifo_cin_PE_3_2_V_V_full_n_pass_0_in = fifo_cin_PE_3_2_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper210_U0_fifo_cin_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper210_U0_fifo_cin_out_V_V_din_pass_0_q0 <= PE_wrapper210_U0_fifo_cin_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper210_U0_fifo_cin_out_V_V_din_pass_0_in = PE_wrapper210_U0_fifo_cin_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper210_U0_fifo_cin_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper210_U0_fifo_cin_out_V_V_write_pass_0_q0 <= PE_wrapper210_U0_fifo_cin_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper210_U0_fifo_cin_out_V_V_write_pass_0_in = PE_wrapper210_U0_fifo_cin_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_cout_drain_IO_L1_out_1_6_V_V_full_n_pass_2_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_cout_drain_IO_L1_out_1_6_V_V_full_n_pass_2_q0 <= fifo_cout_drain_cout_drain_IO_L1_out_1_6_V_V_full_n_pass_2_out;
  end
  assign fifo_cout_drain_cout_drain_IO_L1_out_1_6_V_V_full_n_pass_2_in = fifo_cout_drain_cout_drain_IO_L1_out_1_6_V_V_full_n_pass_2_q0;
  (* dont_touch = "yes" *) reg  ap_done_Boundary_X6Y2_To_X8Y2_q0;
  always @ (posedge ap_clk) begin
    ap_done_Boundary_X6Y2_To_X8Y2_q0 <= ap_done_Boundary_X6Y2_To_X8Y2_out;
  end
  assign ap_done_Boundary_X6Y2_To_X8Y2_in = ap_done_Boundary_X6Y2_To_X8Y2_q0;
  (* dont_touch = "yes" *) reg  ap_start_Boundary_X6Y4_To_X8Y4_q0;
  always @ (posedge ap_clk) begin
    ap_start_Boundary_X6Y4_To_X8Y4_q0 <= ap_start_Boundary_X6Y4_To_X8Y4_out;
  end
  assign ap_start_Boundary_X6Y4_To_X8Y4_in = ap_start_Boundary_X6Y4_To_X8Y4_q0;
  (* dont_touch = "yes" *) reg  ap_rst_n_Boundary_X6Y4_To_X8Y4_q0;
  always @ (posedge ap_clk) begin
    ap_rst_n_Boundary_X6Y4_To_X8Y4_q0 <= ap_rst_n_Boundary_X6Y4_To_X8Y4_out;
  end
  assign ap_rst_n_Boundary_X6Y4_To_X8Y4_in = ap_rst_n_Boundary_X6Y4_To_X8Y4_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper214_U0_fifo_w_out_V_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper214_U0_fifo_w_out_V_V_din_pass_1_q0 <= PE_wrapper214_U0_fifo_w_out_V_V_din_pass_1_out;
  end
  assign PE_wrapper214_U0_fifo_w_out_V_V_din_pass_1_in = PE_wrapper214_U0_fifo_w_out_V_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_5_5_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_5_5_V_V_full_n_pass_0_q0 <= fifo_w_PE_5_5_V_V_full_n_pass_0_out;
  end
  assign fifo_w_PE_5_5_V_V_full_n_pass_0_in = fifo_w_PE_5_5_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper214_U0_fifo_w_out_V_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper214_U0_fifo_w_out_V_V_write_pass_1_q0 <= PE_wrapper214_U0_fifo_w_out_V_V_write_pass_1_out;
  end
  assign PE_wrapper214_U0_fifo_w_out_V_V_write_pass_1_in = PE_wrapper214_U0_fifo_w_out_V_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper202_U0_fifo_w_out_V_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper202_U0_fifo_w_out_V_V_din_pass_1_q0 <= PE_wrapper202_U0_fifo_w_out_V_V_din_pass_1_out;
  end
  assign PE_wrapper202_U0_fifo_w_out_V_V_din_pass_1_in = PE_wrapper202_U0_fifo_w_out_V_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_4_5_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_4_5_V_V_full_n_pass_0_q0 <= fifo_w_PE_4_5_V_V_full_n_pass_0_out;
  end
  assign fifo_w_PE_4_5_V_V_full_n_pass_0_in = fifo_w_PE_4_5_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper202_U0_fifo_w_out_V_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper202_U0_fifo_w_out_V_V_write_pass_1_q0 <= PE_wrapper202_U0_fifo_w_out_V_V_write_pass_1_out;
  end
  assign PE_wrapper202_U0_fifo_w_out_V_V_write_pass_1_in = PE_wrapper202_U0_fifo_w_out_V_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [63:0] kernel0_entry12_U0_cout_V_out_din_pass_3_q0;
  always @ (posedge ap_clk) begin
    kernel0_entry12_U0_cout_V_out_din_pass_3_q0 <= kernel0_entry12_U0_cout_V_out_din_pass_3_out;
  end
  assign kernel0_entry12_U0_cout_V_out_din_pass_3_in = kernel0_entry12_U0_cout_V_out_din_pass_3_q0;
  (* dont_touch = "yes" *) reg  cout_V_c_full_n_pass_2_q0;
  always @ (posedge ap_clk) begin
    cout_V_c_full_n_pass_2_q0 <= cout_V_c_full_n_pass_2_out;
  end
  assign cout_V_c_full_n_pass_2_in = cout_V_c_full_n_pass_2_q0;
  (* dont_touch = "yes" *) reg  kernel0_entry12_U0_cout_V_out_write_pass_3_q0;
  always @ (posedge ap_clk) begin
    kernel0_entry12_U0_cout_V_out_write_pass_3_q0 <= kernel0_entry12_U0_cout_V_out_write_pass_3_out;
  end
  assign kernel0_entry12_U0_cout_V_out_write_pass_3_in = kernel0_entry12_U0_cout_V_out_write_pass_3_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper243_U0_fifo_w_out_V_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper243_U0_fifo_w_out_V_V_din_pass_1_q0 <= PE_wrapper243_U0_fifo_w_out_V_V_din_pass_1_out;
  end
  assign PE_wrapper243_U0_fifo_w_out_V_V_din_pass_1_in = PE_wrapper243_U0_fifo_w_out_V_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_7_10_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_7_10_V_V_full_n_pass_0_q0 <= fifo_w_PE_7_10_V_V_full_n_pass_0_out;
  end
  assign fifo_w_PE_7_10_V_V_full_n_pass_0_in = fifo_w_PE_7_10_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper243_U0_fifo_w_out_V_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper243_U0_fifo_w_out_V_V_write_pass_1_q0 <= PE_wrapper243_U0_fifo_w_out_V_V_write_pass_1_out;
  end
  assign PE_wrapper243_U0_fifo_w_out_V_V_write_pass_1_in = PE_wrapper243_U0_fifo_w_out_V_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [31:0] PE_wrapper243_U0_fifo_cout_drain_out_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper243_U0_fifo_cout_drain_out_V_din_pass_1_q0 <= PE_wrapper243_U0_fifo_cout_drain_out_V_din_pass_1_out;
  end
  assign PE_wrapper243_U0_fifo_cout_drain_out_V_din_pass_1_in = PE_wrapper243_U0_fifo_cout_drain_out_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_PE_7_9_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_PE_7_9_V_full_n_pass_0_q0 <= fifo_cout_drain_PE_7_9_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_PE_7_9_V_full_n_pass_0_in = fifo_cout_drain_PE_7_9_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper243_U0_fifo_cout_drain_out_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper243_U0_fifo_cout_drain_out_V_write_pass_1_q0 <= PE_wrapper243_U0_fifo_cout_drain_out_V_write_pass_1_out;
  end
  assign PE_wrapper243_U0_fifo_cout_drain_out_V_write_pass_1_in = PE_wrapper243_U0_fifo_cout_drain_out_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper243_U0_fifo_cin_out_V_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper243_U0_fifo_cin_out_V_V_din_pass_1_q0 <= PE_wrapper243_U0_fifo_cin_out_V_V_din_pass_1_out;
  end
  assign PE_wrapper243_U0_fifo_cin_out_V_V_din_pass_1_in = PE_wrapper243_U0_fifo_cin_out_V_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_8_9_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_8_9_V_V_full_n_pass_0_q0 <= fifo_cin_PE_8_9_V_V_full_n_pass_0_out;
  end
  assign fifo_cin_PE_8_9_V_V_full_n_pass_0_in = fifo_cin_PE_8_9_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper243_U0_fifo_cin_out_V_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper243_U0_fifo_cin_out_V_V_write_pass_1_q0 <= PE_wrapper243_U0_fifo_cin_out_V_V_write_pass_1_out;
  end
  assign PE_wrapper243_U0_fifo_cin_out_V_V_write_pass_1_in = PE_wrapper243_U0_fifo_cin_out_V_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper191_U0_fifo_cin_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper191_U0_fifo_cin_out_V_V_din_pass_0_q0 <= PE_wrapper191_U0_fifo_cin_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper191_U0_fifo_cin_out_V_V_din_pass_0_in = PE_wrapper191_U0_fifo_cin_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper191_U0_fifo_cin_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper191_U0_fifo_cin_out_V_V_write_pass_0_q0 <= PE_wrapper191_U0_fifo_cin_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper191_U0_fifo_cin_out_V_V_write_pass_0_in = PE_wrapper191_U0_fifo_cin_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [31:0] PE_wrapper191_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper191_U0_fifo_cout_drain_out_V_din_pass_0_q0 <= PE_wrapper191_U0_fifo_cout_drain_out_V_din_pass_0_out;
  end
  assign PE_wrapper191_U0_fifo_cout_drain_out_V_din_pass_0_in = PE_wrapper191_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper191_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper191_U0_fifo_cout_drain_out_V_write_pass_0_q0 <= PE_wrapper191_U0_fifo_cout_drain_out_V_write_pass_0_out;
  end
  assign PE_wrapper191_U0_fifo_cout_drain_out_V_write_pass_0_in = PE_wrapper191_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper192_U0_fifo_cin_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper192_U0_fifo_cin_out_V_V_din_pass_0_q0 <= PE_wrapper192_U0_fifo_cin_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper192_U0_fifo_cin_out_V_V_din_pass_0_in = PE_wrapper192_U0_fifo_cin_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper192_U0_fifo_cin_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper192_U0_fifo_cin_out_V_V_write_pass_0_q0 <= PE_wrapper192_U0_fifo_cin_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper192_U0_fifo_cin_out_V_V_write_pass_0_in = PE_wrapper192_U0_fifo_cin_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [31:0] PE_wrapper192_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper192_U0_fifo_cout_drain_out_V_din_pass_0_q0 <= PE_wrapper192_U0_fifo_cout_drain_out_V_din_pass_0_out;
  end
  assign PE_wrapper192_U0_fifo_cout_drain_out_V_din_pass_0_in = PE_wrapper192_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper192_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper192_U0_fifo_cout_drain_out_V_write_pass_0_q0 <= PE_wrapper192_U0_fifo_cout_drain_out_V_write_pass_0_out;
  end
  assign PE_wrapper192_U0_fifo_cout_drain_out_V_write_pass_0_in = PE_wrapper192_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper192_U0_fifo_w_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper192_U0_fifo_w_out_V_V_din_pass_0_q0 <= PE_wrapper192_U0_fifo_w_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper192_U0_fifo_w_out_V_V_din_pass_0_in = PE_wrapper192_U0_fifo_w_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper192_U0_fifo_w_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper192_U0_fifo_w_out_V_V_write_pass_0_q0 <= PE_wrapper192_U0_fifo_w_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper192_U0_fifo_w_out_V_V_write_pass_0_in = PE_wrapper192_U0_fifo_w_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_3_5_V_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_3_5_V_V_full_n_pass_1_q0 <= fifo_w_PE_3_5_V_V_full_n_pass_1_out;
  end
  assign fifo_w_PE_3_5_V_V_full_n_pass_1_in = fifo_w_PE_3_5_V_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_3_5_V_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_3_5_V_V_full_n_pass_1_q0 <= fifo_cin_PE_3_5_V_V_full_n_pass_1_out;
  end
  assign fifo_cin_PE_3_5_V_V_full_n_pass_1_in = fifo_cin_PE_3_5_V_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_3_6_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_3_6_V_V_full_n_pass_0_q0 <= fifo_cin_PE_3_6_V_V_full_n_pass_0_out;
  end
  assign fifo_cin_PE_3_6_V_V_full_n_pass_0_in = fifo_cin_PE_3_6_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  ap_done_Boundary_X4Y6_To_X6Y6_q0;
  always @ (posedge ap_clk) begin
    ap_done_Boundary_X4Y6_To_X6Y6_q0 <= ap_done_Boundary_X4Y6_To_X6Y6_out;
  end
  assign ap_done_Boundary_X4Y6_To_X6Y6_in = ap_done_Boundary_X4Y6_To_X6Y6_q0;
  (* dont_touch = "yes" *) reg  ap_start_Boundary_X4Y8_To_X6Y8_q0;
  always @ (posedge ap_clk) begin
    ap_start_Boundary_X4Y8_To_X6Y8_q0 <= ap_start_Boundary_X4Y8_To_X6Y8_out;
  end
  assign ap_start_Boundary_X4Y8_To_X6Y8_in = ap_start_Boundary_X4Y8_To_X6Y8_q0;
  (* dont_touch = "yes" *) reg  ap_rst_n_Boundary_X4Y8_To_X6Y8_q0;
  always @ (posedge ap_clk) begin
    ap_rst_n_Boundary_X4Y8_To_X6Y8_q0 <= ap_rst_n_Boundary_X4Y8_To_X6Y8_out;
  end
  assign ap_rst_n_Boundary_X4Y8_To_X6Y8_in = ap_rst_n_Boundary_X4Y8_To_X6Y8_q0;
  (* dont_touch = "yes" *) reg [63:0] cout_drain_IO_L2_out568_U0_fifo_cout_drain_out_V_V_din_pass_2_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L2_out568_U0_fifo_cout_drain_out_V_V_din_pass_2_q0 <= cout_drain_IO_L2_out568_U0_fifo_cout_drain_out_V_V_din_pass_2_out;
  end
  assign cout_drain_IO_L2_out568_U0_fifo_cout_drain_out_V_V_din_pass_2_in = cout_drain_IO_L2_out568_U0_fifo_cout_drain_out_V_V_din_pass_2_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_cout_drain_IO_L2_out_0_V_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_cout_drain_IO_L2_out_0_V_V_full_n_pass_1_q0 <= fifo_cout_drain_cout_drain_IO_L2_out_0_V_V_full_n_pass_1_out;
  end
  assign fifo_cout_drain_cout_drain_IO_L2_out_0_V_V_full_n_pass_1_in = fifo_cout_drain_cout_drain_IO_L2_out_0_V_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg  cout_drain_IO_L2_out568_U0_fifo_cout_drain_out_V_V_write_pass_2_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L2_out568_U0_fifo_cout_drain_out_V_V_write_pass_2_q0 <= cout_drain_IO_L2_out568_U0_fifo_cout_drain_out_V_V_write_pass_2_out;
  end
  assign cout_drain_IO_L2_out568_U0_fifo_cout_drain_out_V_V_write_pass_2_in = cout_drain_IO_L2_out568_U0_fifo_cout_drain_out_V_V_write_pass_2_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_1_4_V_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_1_4_V_V_full_n_pass_1_q0 <= fifo_w_PE_1_4_V_V_full_n_pass_1_out;
  end
  assign fifo_w_PE_1_4_V_V_full_n_pass_1_in = fifo_w_PE_1_4_V_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg [63:0] cout_drain_IO_L2_out564_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L2_out564_U0_fifo_cout_drain_out_V_V_din_pass_0_q0 <= cout_drain_IO_L2_out564_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  end
  assign cout_drain_IO_L2_out564_U0_fifo_cout_drain_out_V_V_din_pass_0_in = cout_drain_IO_L2_out564_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  cout_drain_IO_L2_out564_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L2_out564_U0_fifo_cout_drain_out_V_V_write_pass_0_q0 <= cout_drain_IO_L2_out564_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  end
  assign cout_drain_IO_L2_out564_U0_fifo_cout_drain_out_V_V_write_pass_0_in = cout_drain_IO_L2_out564_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_cin_IO_L2_in_4_V_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_cin_IO_L2_in_4_V_V_full_n_pass_1_q0 <= fifo_cin_cin_IO_L2_in_4_V_V_full_n_pass_1_out;
  end
  assign fifo_cin_cin_IO_L2_in_4_V_V_full_n_pass_1_in = fifo_cin_cin_IO_L2_in_4_V_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper179_U0_fifo_w_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper179_U0_fifo_w_out_V_V_din_pass_0_q0 <= PE_wrapper179_U0_fifo_w_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper179_U0_fifo_w_out_V_V_din_pass_0_in = PE_wrapper179_U0_fifo_w_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper179_U0_fifo_w_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper179_U0_fifo_w_out_V_V_write_pass_0_q0 <= PE_wrapper179_U0_fifo_w_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper179_U0_fifo_w_out_V_V_write_pass_0_in = PE_wrapper179_U0_fifo_w_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] cin_IO_L2_in128_U0_fifo_cin_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    cin_IO_L2_in128_U0_fifo_cin_out_V_V_din_pass_0_q0 <= cin_IO_L2_in128_U0_fifo_cin_out_V_V_din_pass_0_out;
  end
  assign cin_IO_L2_in128_U0_fifo_cin_out_V_V_din_pass_0_in = cin_IO_L2_in128_U0_fifo_cin_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  cin_IO_L2_in128_U0_fifo_cin_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    cin_IO_L2_in128_U0_fifo_cin_out_V_V_write_pass_0_q0 <= cin_IO_L2_in128_U0_fifo_cin_out_V_V_write_pass_0_out;
  end
  assign cin_IO_L2_in128_U0_fifo_cin_out_V_V_write_pass_0_in = cin_IO_L2_in128_U0_fifo_cin_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [31:0] PE_wrapper179_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper179_U0_fifo_cout_drain_out_V_din_pass_0_q0 <= PE_wrapper179_U0_fifo_cout_drain_out_V_din_pass_0_out;
  end
  assign PE_wrapper179_U0_fifo_cout_drain_out_V_din_pass_0_in = PE_wrapper179_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper179_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper179_U0_fifo_cout_drain_out_V_write_pass_0_q0 <= PE_wrapper179_U0_fifo_cout_drain_out_V_write_pass_0_out;
  end
  assign PE_wrapper179_U0_fifo_cout_drain_out_V_write_pass_0_in = PE_wrapper179_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_2_4_V_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_2_4_V_V_full_n_pass_1_q0 <= fifo_w_PE_2_4_V_V_full_n_pass_1_out;
  end
  assign fifo_w_PE_2_4_V_V_full_n_pass_1_in = fifo_w_PE_2_4_V_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_0_4_V_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_0_4_V_V_full_n_pass_1_q0 <= fifo_w_PE_0_4_V_V_full_n_pass_1_out;
  end
  assign fifo_w_PE_0_4_V_V_full_n_pass_1_in = fifo_w_PE_0_4_V_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper190_U0_fifo_cin_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper190_U0_fifo_cin_out_V_V_din_pass_0_q0 <= PE_wrapper190_U0_fifo_cin_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper190_U0_fifo_cin_out_V_V_din_pass_0_in = PE_wrapper190_U0_fifo_cin_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper190_U0_fifo_cin_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper190_U0_fifo_cin_out_V_V_write_pass_0_q0 <= PE_wrapper190_U0_fifo_cin_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper190_U0_fifo_cin_out_V_V_write_pass_0_in = PE_wrapper190_U0_fifo_cin_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper166_U0_fifo_w_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper166_U0_fifo_w_out_V_V_din_pass_0_q0 <= PE_wrapper166_U0_fifo_w_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper166_U0_fifo_w_out_V_V_din_pass_0_in = PE_wrapper166_U0_fifo_w_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper166_U0_fifo_w_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper166_U0_fifo_w_out_V_V_write_pass_0_q0 <= PE_wrapper166_U0_fifo_w_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper166_U0_fifo_w_out_V_V_write_pass_0_in = PE_wrapper166_U0_fifo_w_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper154_U0_fifo_w_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper154_U0_fifo_w_out_V_V_din_pass_0_q0 <= PE_wrapper154_U0_fifo_w_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper154_U0_fifo_w_out_V_V_din_pass_0_in = PE_wrapper154_U0_fifo_w_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper154_U0_fifo_w_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper154_U0_fifo_w_out_V_V_write_pass_0_q0 <= PE_wrapper154_U0_fifo_w_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper154_U0_fifo_w_out_V_V_write_pass_0_in = PE_wrapper154_U0_fifo_w_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_cout_drain_IO_L2_out_5_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_cout_drain_IO_L2_out_5_V_V_full_n_pass_0_q0 <= fifo_cout_drain_cout_drain_IO_L2_out_5_V_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_cout_drain_IO_L2_out_5_V_V_full_n_pass_0_in = fifo_cout_drain_cout_drain_IO_L2_out_5_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper190_U0_fifo_w_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper190_U0_fifo_w_out_V_V_din_pass_0_q0 <= PE_wrapper190_U0_fifo_w_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper190_U0_fifo_w_out_V_V_din_pass_0_in = PE_wrapper190_U0_fifo_w_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper190_U0_fifo_w_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper190_U0_fifo_w_out_V_V_write_pass_0_q0 <= PE_wrapper190_U0_fifo_w_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper190_U0_fifo_w_out_V_V_write_pass_0_in = PE_wrapper190_U0_fifo_w_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper179_U0_fifo_cin_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper179_U0_fifo_cin_out_V_V_din_pass_0_q0 <= PE_wrapper179_U0_fifo_cin_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper179_U0_fifo_cin_out_V_V_din_pass_0_in = PE_wrapper179_U0_fifo_cin_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper179_U0_fifo_cin_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper179_U0_fifo_cin_out_V_V_write_pass_0_q0 <= PE_wrapper179_U0_fifo_cin_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper179_U0_fifo_cin_out_V_V_write_pass_0_in = PE_wrapper179_U0_fifo_cin_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_PE_4_4_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_PE_4_4_V_full_n_pass_0_q0 <= fifo_cout_drain_PE_4_4_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_PE_4_4_V_full_n_pass_0_in = fifo_cout_drain_PE_4_4_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_3_4_V_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_3_4_V_V_full_n_pass_1_q0 <= fifo_w_PE_3_4_V_V_full_n_pass_1_out;
  end
  assign fifo_w_PE_3_4_V_V_full_n_pass_1_in = fifo_w_PE_3_4_V_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_2_5_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_2_5_V_V_full_n_pass_0_q0 <= fifo_cin_PE_2_5_V_V_full_n_pass_0_out;
  end
  assign fifo_cin_PE_2_5_V_V_full_n_pass_0_in = fifo_cin_PE_2_5_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_cout_drain_IO_L1_out_4_5_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_cout_drain_IO_L1_out_4_5_V_V_full_n_pass_0_q0 <= fifo_cout_drain_cout_drain_IO_L1_out_4_5_V_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_cout_drain_IO_L1_out_4_5_V_V_full_n_pass_0_in = fifo_cout_drain_cout_drain_IO_L1_out_4_5_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  ap_done_Boundary_X6Y4_To_X8Y4_q0;
  always @ (posedge ap_clk) begin
    ap_done_Boundary_X6Y4_To_X8Y4_q0 <= ap_done_Boundary_X6Y4_To_X8Y4_out;
  end
  assign ap_done_Boundary_X6Y4_To_X8Y4_in = ap_done_Boundary_X6Y4_To_X8Y4_q0;
  (* dont_touch = "yes" *) reg  ap_start_Boundary_X6Y6_To_X8Y6_q0;
  always @ (posedge ap_clk) begin
    ap_start_Boundary_X6Y6_To_X8Y6_q0 <= ap_start_Boundary_X6Y6_To_X8Y6_out;
  end
  assign ap_start_Boundary_X6Y6_To_X8Y6_in = ap_start_Boundary_X6Y6_To_X8Y6_q0;
  (* dont_touch = "yes" *) reg  ap_rst_n_Boundary_X6Y6_To_X8Y6_q0;
  always @ (posedge ap_clk) begin
    ap_rst_n_Boundary_X6Y6_To_X8Y6_q0 <= ap_rst_n_Boundary_X6Y6_To_X8Y6_out;
  end
  assign ap_rst_n_Boundary_X6Y6_To_X8Y6_in = ap_rst_n_Boundary_X6Y6_To_X8Y6_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper192_U0_fifo_w_out_V_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper192_U0_fifo_w_out_V_V_din_pass_1_q0 <= PE_wrapper192_U0_fifo_w_out_V_V_din_pass_1_out;
  end
  assign PE_wrapper192_U0_fifo_w_out_V_V_din_pass_1_in = PE_wrapper192_U0_fifo_w_out_V_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_3_7_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_3_7_V_V_full_n_pass_0_q0 <= fifo_w_PE_3_7_V_V_full_n_pass_0_out;
  end
  assign fifo_w_PE_3_7_V_V_full_n_pass_0_in = fifo_w_PE_3_7_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper192_U0_fifo_w_out_V_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper192_U0_fifo_w_out_V_V_write_pass_1_q0 <= PE_wrapper192_U0_fifo_w_out_V_V_write_pass_1_out;
  end
  assign PE_wrapper192_U0_fifo_w_out_V_V_write_pass_1_in = PE_wrapper192_U0_fifo_w_out_V_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [63:0] cout_drain_IO_L2_out568_U0_fifo_cout_drain_out_V_V_din_pass_3_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L2_out568_U0_fifo_cout_drain_out_V_V_din_pass_3_q0 <= cout_drain_IO_L2_out568_U0_fifo_cout_drain_out_V_V_din_pass_3_out;
  end
  assign cout_drain_IO_L2_out568_U0_fifo_cout_drain_out_V_V_din_pass_3_in = cout_drain_IO_L2_out568_U0_fifo_cout_drain_out_V_V_din_pass_3_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_cout_drain_IO_L2_out_0_V_V_full_n_pass_2_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_cout_drain_IO_L2_out_0_V_V_full_n_pass_2_q0 <= fifo_cout_drain_cout_drain_IO_L2_out_0_V_V_full_n_pass_2_out;
  end
  assign fifo_cout_drain_cout_drain_IO_L2_out_0_V_V_full_n_pass_2_in = fifo_cout_drain_cout_drain_IO_L2_out_0_V_V_full_n_pass_2_q0;
  (* dont_touch = "yes" *) reg  cout_drain_IO_L2_out568_U0_fifo_cout_drain_out_V_V_write_pass_3_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L2_out568_U0_fifo_cout_drain_out_V_V_write_pass_3_q0 <= cout_drain_IO_L2_out568_U0_fifo_cout_drain_out_V_V_write_pass_3_out;
  end
  assign cout_drain_IO_L2_out568_U0_fifo_cout_drain_out_V_V_write_pass_3_in = cout_drain_IO_L2_out568_U0_fifo_cout_drain_out_V_V_write_pass_3_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper168_U0_fifo_w_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper168_U0_fifo_w_out_V_V_din_pass_0_q0 <= PE_wrapper168_U0_fifo_w_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper168_U0_fifo_w_out_V_V_din_pass_0_in = PE_wrapper168_U0_fifo_w_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper168_U0_fifo_w_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper168_U0_fifo_w_out_V_V_write_pass_0_q0 <= PE_wrapper168_U0_fifo_w_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper168_U0_fifo_w_out_V_V_write_pass_0_in = PE_wrapper168_U0_fifo_w_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_2_6_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_2_6_V_V_full_n_pass_0_q0 <= fifo_w_PE_2_6_V_V_full_n_pass_0_out;
  end
  assign fifo_w_PE_2_6_V_V_full_n_pass_0_in = fifo_w_PE_2_6_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_cin_IO_L2_in_5_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_cin_IO_L2_in_5_V_V_full_n_pass_0_q0 <= fifo_cin_cin_IO_L2_in_5_V_V_full_n_pass_0_out;
  end
  assign fifo_cin_cin_IO_L2_in_5_V_V_full_n_pass_0_in = fifo_cin_cin_IO_L2_in_5_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_cout_drain_IO_L2_out_7_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_cout_drain_IO_L2_out_7_V_V_full_n_pass_0_q0 <= fifo_cout_drain_cout_drain_IO_L2_out_7_V_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_cout_drain_IO_L2_out_7_V_V_full_n_pass_0_in = fifo_cout_drain_cout_drain_IO_L2_out_7_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_7_9_V_V_full_n_pass_2_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_7_9_V_V_full_n_pass_2_q0 <= fifo_w_PE_7_9_V_V_full_n_pass_2_out;
  end
  assign fifo_w_PE_7_9_V_V_full_n_pass_2_in = fifo_w_PE_7_9_V_V_full_n_pass_2_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_PE_2_5_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_PE_2_5_V_full_n_pass_0_q0 <= fifo_cout_drain_PE_2_5_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_PE_2_5_V_full_n_pass_0_in = fifo_cout_drain_PE_2_5_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] cin_IO_L2_in130_U0_fifo_cin_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    cin_IO_L2_in130_U0_fifo_cin_out_V_V_din_pass_0_q0 <= cin_IO_L2_in130_U0_fifo_cin_out_V_V_din_pass_0_out;
  end
  assign cin_IO_L2_in130_U0_fifo_cin_out_V_V_din_pass_0_in = cin_IO_L2_in130_U0_fifo_cin_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  cin_IO_L2_in130_U0_fifo_cin_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    cin_IO_L2_in130_U0_fifo_cin_out_V_V_write_pass_0_q0 <= cin_IO_L2_in130_U0_fifo_cin_out_V_V_write_pass_0_out;
  end
  assign cin_IO_L2_in130_U0_fifo_cin_out_V_V_write_pass_0_in = cin_IO_L2_in130_U0_fifo_cin_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_1_5_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_1_5_V_V_full_n_pass_0_q0 <= fifo_w_PE_1_5_V_V_full_n_pass_0_out;
  end
  assign fifo_w_PE_1_5_V_V_full_n_pass_0_in = fifo_w_PE_1_5_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper243_U0_fifo_w_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper243_U0_fifo_w_out_V_V_din_pass_0_q0 <= PE_wrapper243_U0_fifo_w_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper243_U0_fifo_w_out_V_V_din_pass_0_in = PE_wrapper243_U0_fifo_w_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper243_U0_fifo_w_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper243_U0_fifo_w_out_V_V_write_pass_0_q0 <= PE_wrapper243_U0_fifo_w_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper243_U0_fifo_w_out_V_V_write_pass_0_in = PE_wrapper243_U0_fifo_w_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [31:0] PE_wrapper243_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper243_U0_fifo_cout_drain_out_V_din_pass_0_q0 <= PE_wrapper243_U0_fifo_cout_drain_out_V_din_pass_0_out;
  end
  assign PE_wrapper243_U0_fifo_cout_drain_out_V_din_pass_0_in = PE_wrapper243_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper243_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper243_U0_fifo_cout_drain_out_V_write_pass_0_q0 <= PE_wrapper243_U0_fifo_cout_drain_out_V_write_pass_0_out;
  end
  assign PE_wrapper243_U0_fifo_cout_drain_out_V_write_pass_0_in = PE_wrapper243_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper243_U0_fifo_cin_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper243_U0_fifo_cin_out_V_V_din_pass_0_q0 <= PE_wrapper243_U0_fifo_cin_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper243_U0_fifo_cin_out_V_V_din_pass_0_in = PE_wrapper243_U0_fifo_cin_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper243_U0_fifo_cin_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper243_U0_fifo_cin_out_V_V_write_pass_0_q0 <= PE_wrapper243_U0_fifo_cin_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper243_U0_fifo_cin_out_V_V_write_pass_0_in = PE_wrapper243_U0_fifo_cin_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_0_5_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_0_5_V_V_full_n_pass_0_q0 <= fifo_w_PE_0_5_V_V_full_n_pass_0_out;
  end
  assign fifo_w_PE_0_5_V_V_full_n_pass_0_in = fifo_w_PE_0_5_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper156_U0_fifo_w_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper156_U0_fifo_w_out_V_V_din_pass_0_q0 <= PE_wrapper156_U0_fifo_w_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper156_U0_fifo_w_out_V_V_din_pass_0_in = PE_wrapper156_U0_fifo_w_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper156_U0_fifo_w_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper156_U0_fifo_w_out_V_V_write_pass_0_q0 <= PE_wrapper156_U0_fifo_w_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper156_U0_fifo_w_out_V_V_write_pass_0_in = PE_wrapper156_U0_fifo_w_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper180_U0_fifo_cin_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper180_U0_fifo_cin_out_V_V_din_pass_0_q0 <= PE_wrapper180_U0_fifo_cin_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper180_U0_fifo_cin_out_V_V_din_pass_0_in = PE_wrapper180_U0_fifo_cin_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper180_U0_fifo_cin_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper180_U0_fifo_cin_out_V_V_write_pass_0_q0 <= PE_wrapper180_U0_fifo_cin_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper180_U0_fifo_cin_out_V_V_write_pass_0_in = PE_wrapper180_U0_fifo_cin_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [63:0] cout_drain_IO_L2_out563_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L2_out563_U0_fifo_cout_drain_out_V_V_din_pass_0_q0 <= cout_drain_IO_L2_out563_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  end
  assign cout_drain_IO_L2_out563_U0_fifo_cout_drain_out_V_V_din_pass_0_in = cout_drain_IO_L2_out563_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  cout_drain_IO_L2_out563_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L2_out563_U0_fifo_cout_drain_out_V_V_write_pass_0_q0 <= cout_drain_IO_L2_out563_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  end
  assign cout_drain_IO_L2_out563_U0_fifo_cout_drain_out_V_V_write_pass_0_in = cout_drain_IO_L2_out563_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_PE_3_5_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_PE_3_5_V_full_n_pass_0_q0 <= fifo_cout_drain_PE_3_5_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_PE_3_5_V_full_n_pass_0_in = fifo_cout_drain_PE_3_5_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_cout_drain_IO_L1_out_6_4_V_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_cout_drain_IO_L1_out_6_4_V_V_full_n_pass_1_q0 <= fifo_cout_drain_cout_drain_IO_L1_out_6_4_V_V_full_n_pass_1_out;
  end
  assign fifo_cout_drain_cout_drain_IO_L1_out_6_4_V_V_full_n_pass_1_in = fifo_cout_drain_cout_drain_IO_L1_out_6_4_V_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_cout_drain_IO_L1_out_5_4_V_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_cout_drain_IO_L1_out_5_4_V_V_full_n_pass_1_q0 <= fifo_cout_drain_cout_drain_IO_L1_out_5_4_V_V_full_n_pass_1_out;
  end
  assign fifo_cout_drain_cout_drain_IO_L1_out_5_4_V_V_full_n_pass_1_in = fifo_cout_drain_cout_drain_IO_L1_out_5_4_V_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper180_U0_fifo_w_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper180_U0_fifo_w_out_V_V_din_pass_0_q0 <= PE_wrapper180_U0_fifo_w_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper180_U0_fifo_w_out_V_V_din_pass_0_in = PE_wrapper180_U0_fifo_w_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper180_U0_fifo_w_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper180_U0_fifo_w_out_V_V_write_pass_0_q0 <= PE_wrapper180_U0_fifo_w_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper180_U0_fifo_w_out_V_V_write_pass_0_in = PE_wrapper180_U0_fifo_w_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper167_U0_fifo_cin_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper167_U0_fifo_cin_out_V_V_din_pass_0_q0 <= PE_wrapper167_U0_fifo_cin_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper167_U0_fifo_cin_out_V_V_din_pass_0_in = PE_wrapper167_U0_fifo_cin_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper167_U0_fifo_cin_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper167_U0_fifo_cin_out_V_V_write_pass_0_q0 <= PE_wrapper167_U0_fifo_cin_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper167_U0_fifo_cin_out_V_V_write_pass_0_in = PE_wrapper167_U0_fifo_cin_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_PE_3_6_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_PE_3_6_V_full_n_pass_0_q0 <= fifo_cout_drain_PE_3_6_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_PE_3_6_V_full_n_pass_0_in = fifo_cout_drain_PE_3_6_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_7_9_V_V_full_n_pass_4_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_7_9_V_V_full_n_pass_4_q0 <= fifo_cin_PE_7_9_V_V_full_n_pass_4_out;
  end
  assign fifo_cin_PE_7_9_V_V_full_n_pass_4_in = fifo_cin_PE_7_9_V_V_full_n_pass_4_q0;
  (* dont_touch = "yes" *) reg  ap_done_Boundary_X6Y6_To_X8Y6_q0;
  always @ (posedge ap_clk) begin
    ap_done_Boundary_X6Y6_To_X8Y6_q0 <= ap_done_Boundary_X6Y6_To_X8Y6_out;
  end
  assign ap_done_Boundary_X6Y6_To_X8Y6_in = ap_done_Boundary_X6Y6_To_X8Y6_q0;
  (* dont_touch = "yes" *) reg  ap_start_Boundary_X6Y8_To_X8Y8_q0;
  always @ (posedge ap_clk) begin
    ap_start_Boundary_X6Y8_To_X8Y8_q0 <= ap_start_Boundary_X6Y8_To_X8Y8_out;
  end
  assign ap_start_Boundary_X6Y8_To_X8Y8_in = ap_start_Boundary_X6Y8_To_X8Y8_q0;
  (* dont_touch = "yes" *) reg  ap_rst_n_Boundary_X6Y8_To_X8Y8_q0;
  always @ (posedge ap_clk) begin
    ap_rst_n_Boundary_X6Y8_To_X8Y8_q0 <= ap_rst_n_Boundary_X6Y8_To_X8Y8_out;
  end
  assign ap_rst_n_Boundary_X6Y8_To_X8Y8_in = ap_rst_n_Boundary_X6Y8_To_X8Y8_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper251_U0_fifo_w_out_V_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper251_U0_fifo_w_out_V_V_din_pass_1_q0 <= PE_wrapper251_U0_fifo_w_out_V_V_din_pass_1_out;
  end
  assign PE_wrapper251_U0_fifo_w_out_V_V_din_pass_1_in = PE_wrapper251_U0_fifo_w_out_V_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_8_6_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_8_6_V_V_full_n_pass_0_q0 <= fifo_w_PE_8_6_V_V_full_n_pass_0_out;
  end
  assign fifo_w_PE_8_6_V_V_full_n_pass_0_in = fifo_w_PE_8_6_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper251_U0_fifo_w_out_V_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper251_U0_fifo_w_out_V_V_write_pass_1_q0 <= PE_wrapper251_U0_fifo_w_out_V_V_write_pass_1_out;
  end
  assign PE_wrapper251_U0_fifo_w_out_V_V_write_pass_1_in = PE_wrapper251_U0_fifo_w_out_V_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper239_U0_fifo_w_out_V_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper239_U0_fifo_w_out_V_V_din_pass_1_q0 <= PE_wrapper239_U0_fifo_w_out_V_V_din_pass_1_out;
  end
  assign PE_wrapper239_U0_fifo_w_out_V_V_din_pass_1_in = PE_wrapper239_U0_fifo_w_out_V_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_7_6_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_7_6_V_V_full_n_pass_0_q0 <= fifo_w_PE_7_6_V_V_full_n_pass_0_out;
  end
  assign fifo_w_PE_7_6_V_V_full_n_pass_0_in = fifo_w_PE_7_6_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper239_U0_fifo_w_out_V_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper239_U0_fifo_w_out_V_V_write_pass_1_q0 <= PE_wrapper239_U0_fifo_w_out_V_V_write_pass_1_out;
  end
  assign PE_wrapper239_U0_fifo_w_out_V_V_write_pass_1_in = PE_wrapper239_U0_fifo_w_out_V_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [63:0] cout_drain_IO_L1_out_wrapper469_U0_fifo_cout_drain_out_V_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper469_U0_fifo_cout_drain_out_V_V_din_pass_1_q0 <= cout_drain_IO_L1_out_wrapper469_U0_fifo_cout_drain_out_V_V_din_pass_1_out;
  end
  assign cout_drain_IO_L1_out_wrapper469_U0_fifo_cout_drain_out_V_V_din_pass_1_in = cout_drain_IO_L1_out_wrapper469_U0_fifo_cout_drain_out_V_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_cout_drain_IO_L1_out_6_9_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_cout_drain_IO_L1_out_6_9_V_V_full_n_pass_0_q0 <= fifo_cout_drain_cout_drain_IO_L1_out_6_9_V_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_cout_drain_IO_L1_out_6_9_V_V_full_n_pass_0_in = fifo_cout_drain_cout_drain_IO_L1_out_6_9_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  cout_drain_IO_L1_out_wrapper469_U0_fifo_cout_drain_out_V_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper469_U0_fifo_cout_drain_out_V_V_write_pass_1_q0 <= cout_drain_IO_L1_out_wrapper469_U0_fifo_cout_drain_out_V_V_write_pass_1_out;
  end
  assign cout_drain_IO_L1_out_wrapper469_U0_fifo_cout_drain_out_V_V_write_pass_1_in = cout_drain_IO_L1_out_wrapper469_U0_fifo_cout_drain_out_V_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [63:0] kernel0_entry12_U0_cout_V_out_din_pass_4_q0;
  always @ (posedge ap_clk) begin
    kernel0_entry12_U0_cout_V_out_din_pass_4_q0 <= kernel0_entry12_U0_cout_V_out_din_pass_4_out;
  end
  assign kernel0_entry12_U0_cout_V_out_din_pass_4_in = kernel0_entry12_U0_cout_V_out_din_pass_4_q0;
  (* dont_touch = "yes" *) reg  cout_V_c_full_n_pass_3_q0;
  always @ (posedge ap_clk) begin
    cout_V_c_full_n_pass_3_q0 <= cout_V_c_full_n_pass_3_out;
  end
  assign cout_V_c_full_n_pass_3_in = cout_V_c_full_n_pass_3_q0;
  (* dont_touch = "yes" *) reg  kernel0_entry12_U0_cout_V_out_write_pass_4_q0;
  always @ (posedge ap_clk) begin
    kernel0_entry12_U0_cout_V_out_write_pass_4_q0 <= kernel0_entry12_U0_cout_V_out_write_pass_4_out;
  end
  assign kernel0_entry12_U0_cout_V_out_write_pass_4_in = kernel0_entry12_U0_cout_V_out_write_pass_4_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper243_U0_fifo_w_out_V_V_din_pass_2_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper243_U0_fifo_w_out_V_V_din_pass_2_q0 <= PE_wrapper243_U0_fifo_w_out_V_V_din_pass_2_out;
  end
  assign PE_wrapper243_U0_fifo_w_out_V_V_din_pass_2_in = PE_wrapper243_U0_fifo_w_out_V_V_din_pass_2_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_7_10_V_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_7_10_V_V_full_n_pass_1_q0 <= fifo_w_PE_7_10_V_V_full_n_pass_1_out;
  end
  assign fifo_w_PE_7_10_V_V_full_n_pass_1_in = fifo_w_PE_7_10_V_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper243_U0_fifo_w_out_V_V_write_pass_2_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper243_U0_fifo_w_out_V_V_write_pass_2_q0 <= PE_wrapper243_U0_fifo_w_out_V_V_write_pass_2_out;
  end
  assign PE_wrapper243_U0_fifo_w_out_V_V_write_pass_2_in = PE_wrapper243_U0_fifo_w_out_V_V_write_pass_2_q0;
  (* dont_touch = "yes" *) reg [31:0] PE_wrapper243_U0_fifo_cout_drain_out_V_din_pass_2_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper243_U0_fifo_cout_drain_out_V_din_pass_2_q0 <= PE_wrapper243_U0_fifo_cout_drain_out_V_din_pass_2_out;
  end
  assign PE_wrapper243_U0_fifo_cout_drain_out_V_din_pass_2_in = PE_wrapper243_U0_fifo_cout_drain_out_V_din_pass_2_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_PE_7_9_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_PE_7_9_V_full_n_pass_1_q0 <= fifo_cout_drain_PE_7_9_V_full_n_pass_1_out;
  end
  assign fifo_cout_drain_PE_7_9_V_full_n_pass_1_in = fifo_cout_drain_PE_7_9_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper243_U0_fifo_cout_drain_out_V_write_pass_2_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper243_U0_fifo_cout_drain_out_V_write_pass_2_q0 <= PE_wrapper243_U0_fifo_cout_drain_out_V_write_pass_2_out;
  end
  assign PE_wrapper243_U0_fifo_cout_drain_out_V_write_pass_2_in = PE_wrapper243_U0_fifo_cout_drain_out_V_write_pass_2_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper243_U0_fifo_cin_out_V_V_din_pass_2_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper243_U0_fifo_cin_out_V_V_din_pass_2_q0 <= PE_wrapper243_U0_fifo_cin_out_V_V_din_pass_2_out;
  end
  assign PE_wrapper243_U0_fifo_cin_out_V_V_din_pass_2_in = PE_wrapper243_U0_fifo_cin_out_V_V_din_pass_2_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_8_9_V_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_8_9_V_V_full_n_pass_1_q0 <= fifo_cin_PE_8_9_V_V_full_n_pass_1_out;
  end
  assign fifo_cin_PE_8_9_V_V_full_n_pass_1_in = fifo_cin_PE_8_9_V_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper243_U0_fifo_cin_out_V_V_write_pass_2_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper243_U0_fifo_cin_out_V_V_write_pass_2_q0 <= PE_wrapper243_U0_fifo_cin_out_V_V_write_pass_2_out;
  end
  assign PE_wrapper243_U0_fifo_cin_out_V_V_write_pass_2_in = PE_wrapper243_U0_fifo_cin_out_V_V_write_pass_2_q0;
  (* dont_touch = "yes" *) reg [63:0] cout_drain_IO_L3_out_U0_fifo_cout_drain_out_V_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L3_out_U0_fifo_cout_drain_out_V_V_din_pass_1_q0 <= cout_drain_IO_L3_out_U0_fifo_cout_drain_out_V_V_din_pass_1_out;
  end
  assign cout_drain_IO_L3_out_U0_fifo_cout_drain_out_V_V_din_pass_1_in = cout_drain_IO_L3_out_U0_fifo_cout_drain_out_V_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_cout_drain_IO_L3_out_serialize_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_cout_drain_IO_L3_out_serialize_V_V_full_n_pass_0_q0 <= fifo_cout_drain_cout_drain_IO_L3_out_serialize_V_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_cout_drain_IO_L3_out_serialize_V_V_full_n_pass_0_in = fifo_cout_drain_cout_drain_IO_L3_out_serialize_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  cout_drain_IO_L3_out_U0_fifo_cout_drain_out_V_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L3_out_U0_fifo_cout_drain_out_V_V_write_pass_1_q0 <= cout_drain_IO_L3_out_U0_fifo_cout_drain_out_V_V_write_pass_1_out;
  end
  assign cout_drain_IO_L3_out_U0_fifo_cout_drain_out_V_V_write_pass_1_in = cout_drain_IO_L3_out_U0_fifo_cout_drain_out_V_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_4_6_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_4_6_V_V_full_n_pass_0_q0 <= fifo_cin_PE_4_6_V_V_full_n_pass_0_out;
  end
  assign fifo_cin_PE_4_6_V_V_full_n_pass_0_in = fifo_cin_PE_4_6_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_cout_drain_IO_L1_out_6_7_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_cout_drain_IO_L1_out_6_7_V_V_full_n_pass_0_q0 <= fifo_cout_drain_cout_drain_IO_L1_out_6_7_V_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_cout_drain_IO_L1_out_6_7_V_V_full_n_pass_0_in = fifo_cout_drain_cout_drain_IO_L1_out_6_7_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_5_5_V_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_5_5_V_V_full_n_pass_1_q0 <= fifo_w_PE_5_5_V_V_full_n_pass_1_out;
  end
  assign fifo_w_PE_5_5_V_V_full_n_pass_1_in = fifo_w_PE_5_5_V_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg [63:0] cout_drain_IO_L1_out_wrapper490_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper490_U0_fifo_cout_drain_out_V_V_din_pass_0_q0 <= cout_drain_IO_L1_out_wrapper490_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper490_U0_fifo_cout_drain_out_V_V_din_pass_0_in = cout_drain_IO_L1_out_wrapper490_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  cout_drain_IO_L1_out_wrapper490_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper490_U0_fifo_cout_drain_out_V_V_write_pass_0_q0 <= cout_drain_IO_L1_out_wrapper490_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper490_U0_fifo_cout_drain_out_V_V_write_pass_0_in = cout_drain_IO_L1_out_wrapper490_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_5_7_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_5_7_V_V_full_n_pass_0_q0 <= fifo_cin_PE_5_7_V_V_full_n_pass_0_out;
  end
  assign fifo_cin_PE_5_7_V_V_full_n_pass_0_in = fifo_cin_PE_5_7_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper217_U0_fifo_w_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper217_U0_fifo_w_out_V_V_din_pass_0_q0 <= PE_wrapper217_U0_fifo_w_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper217_U0_fifo_w_out_V_V_din_pass_0_in = PE_wrapper217_U0_fifo_w_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper217_U0_fifo_w_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper217_U0_fifo_w_out_V_V_write_pass_0_q0 <= PE_wrapper217_U0_fifo_w_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper217_U0_fifo_w_out_V_V_write_pass_0_in = PE_wrapper217_U0_fifo_w_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper215_U0_fifo_cin_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper215_U0_fifo_cin_out_V_V_din_pass_0_q0 <= PE_wrapper215_U0_fifo_cin_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper215_U0_fifo_cin_out_V_V_din_pass_0_in = PE_wrapper215_U0_fifo_cin_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper215_U0_fifo_cin_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper215_U0_fifo_cin_out_V_V_write_pass_0_q0 <= PE_wrapper215_U0_fifo_cin_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper215_U0_fifo_cin_out_V_V_write_pass_0_in = PE_wrapper215_U0_fifo_cin_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_6_6_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_6_6_V_V_full_n_pass_0_q0 <= fifo_w_PE_6_6_V_V_full_n_pass_0_out;
  end
  assign fifo_w_PE_6_6_V_V_full_n_pass_0_in = fifo_w_PE_6_6_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper228_U0_fifo_cin_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper228_U0_fifo_cin_out_V_V_din_pass_0_q0 <= PE_wrapper228_U0_fifo_cin_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper228_U0_fifo_cin_out_V_V_din_pass_0_in = PE_wrapper228_U0_fifo_cin_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper228_U0_fifo_cin_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper228_U0_fifo_cin_out_V_V_write_pass_0_q0 <= PE_wrapper228_U0_fifo_cin_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper228_U0_fifo_cin_out_V_V_write_pass_0_in = PE_wrapper228_U0_fifo_cin_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [63:0] cout_drain_IO_L1_out_wrapper474_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper474_U0_fifo_cout_drain_out_V_V_din_pass_0_q0 <= cout_drain_IO_L1_out_wrapper474_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper474_U0_fifo_cout_drain_out_V_V_din_pass_0_in = cout_drain_IO_L1_out_wrapper474_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  cout_drain_IO_L1_out_wrapper474_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper474_U0_fifo_cout_drain_out_V_V_write_pass_0_q0 <= cout_drain_IO_L1_out_wrapper474_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper474_U0_fifo_cout_drain_out_V_V_write_pass_0_in = cout_drain_IO_L1_out_wrapper474_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [63:0] cout_drain_IO_L1_out_wrapper458_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper458_U0_fifo_cout_drain_out_V_V_din_pass_0_q0 <= cout_drain_IO_L1_out_wrapper458_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper458_U0_fifo_cout_drain_out_V_V_din_pass_0_in = cout_drain_IO_L1_out_wrapper458_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  cout_drain_IO_L1_out_wrapper458_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper458_U0_fifo_cout_drain_out_V_V_write_pass_0_q0 <= cout_drain_IO_L1_out_wrapper458_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper458_U0_fifo_cout_drain_out_V_V_write_pass_0_in = cout_drain_IO_L1_out_wrapper458_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper229_U0_fifo_w_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper229_U0_fifo_w_out_V_V_din_pass_0_q0 <= PE_wrapper229_U0_fifo_w_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper229_U0_fifo_w_out_V_V_din_pass_0_in = PE_wrapper229_U0_fifo_w_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper229_U0_fifo_w_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper229_U0_fifo_w_out_V_V_write_pass_0_q0 <= PE_wrapper229_U0_fifo_w_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper229_U0_fifo_w_out_V_V_write_pass_0_in = PE_wrapper229_U0_fifo_w_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_4_5_V_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_4_5_V_V_full_n_pass_1_q0 <= fifo_w_PE_4_5_V_V_full_n_pass_1_out;
  end
  assign fifo_w_PE_4_5_V_V_full_n_pass_1_in = fifo_w_PE_4_5_V_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_cout_drain_IO_L1_out_5_6_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_cout_drain_IO_L1_out_5_6_V_V_full_n_pass_0_q0 <= fifo_cout_drain_cout_drain_IO_L1_out_5_6_V_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_cout_drain_IO_L1_out_5_6_V_V_full_n_pass_0_in = fifo_cout_drain_cout_drain_IO_L1_out_5_6_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper229_U0_fifo_cin_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper229_U0_fifo_cin_out_V_V_din_pass_0_q0 <= PE_wrapper229_U0_fifo_cin_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper229_U0_fifo_cin_out_V_V_din_pass_0_in = PE_wrapper229_U0_fifo_cin_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper229_U0_fifo_cin_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper229_U0_fifo_cin_out_V_V_write_pass_0_q0 <= PE_wrapper229_U0_fifo_cin_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper229_U0_fifo_cin_out_V_V_write_pass_0_in = PE_wrapper229_U0_fifo_cin_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_4_5_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_4_5_V_V_full_n_pass_0_q0 <= fifo_cin_PE_4_5_V_V_full_n_pass_0_out;
  end
  assign fifo_cin_PE_4_5_V_V_full_n_pass_0_in = fifo_cin_PE_4_5_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_PE_4_7_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_PE_4_7_V_full_n_pass_0_q0 <= fifo_cout_drain_PE_4_7_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_PE_4_7_V_full_n_pass_0_in = fifo_cout_drain_PE_4_7_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper204_U0_fifo_w_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper204_U0_fifo_w_out_V_V_din_pass_0_q0 <= PE_wrapper204_U0_fifo_w_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper204_U0_fifo_w_out_V_V_din_pass_0_in = PE_wrapper204_U0_fifo_w_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper204_U0_fifo_w_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper204_U0_fifo_w_out_V_V_write_pass_0_q0 <= PE_wrapper204_U0_fifo_w_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper204_U0_fifo_w_out_V_V_write_pass_0_in = PE_wrapper204_U0_fifo_w_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_cout_drain_IO_L1_out_7_7_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_cout_drain_IO_L1_out_7_7_V_V_full_n_pass_0_q0 <= fifo_cout_drain_cout_drain_IO_L1_out_7_7_V_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_cout_drain_IO_L1_out_7_7_V_V_full_n_pass_0_in = fifo_cout_drain_cout_drain_IO_L1_out_7_7_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  ap_done_Boundary_X4Y8_To_X6Y8_q0;
  always @ (posedge ap_clk) begin
    ap_done_Boundary_X4Y8_To_X6Y8_q0 <= ap_done_Boundary_X4Y8_To_X6Y8_out;
  end
  assign ap_done_Boundary_X4Y8_To_X6Y8_in = ap_done_Boundary_X4Y8_To_X6Y8_q0;
  (* dont_touch = "yes" *) reg  ap_start_Boundary_X4Y10_To_X6Y10_q0;
  always @ (posedge ap_clk) begin
    ap_start_Boundary_X4Y10_To_X6Y10_q0 <= ap_start_Boundary_X4Y10_To_X6Y10_out;
  end
  assign ap_start_Boundary_X4Y10_To_X6Y10_in = ap_start_Boundary_X4Y10_To_X6Y10_q0;
  (* dont_touch = "yes" *) reg  ap_rst_n_Boundary_X4Y10_To_X6Y10_q0;
  always @ (posedge ap_clk) begin
    ap_rst_n_Boundary_X4Y10_To_X6Y10_q0 <= ap_rst_n_Boundary_X4Y10_To_X6Y10_out;
  end
  assign ap_rst_n_Boundary_X4Y10_To_X6Y10_in = ap_rst_n_Boundary_X4Y10_To_X6Y10_q0;
  (* dont_touch = "yes" *) reg [63:0] kernel0_entry12_U0_cout_V_out_din_pass_5_q0;
  always @ (posedge ap_clk) begin
    kernel0_entry12_U0_cout_V_out_din_pass_5_q0 <= kernel0_entry12_U0_cout_V_out_din_pass_5_out;
  end
  assign kernel0_entry12_U0_cout_V_out_din_pass_5_in = kernel0_entry12_U0_cout_V_out_din_pass_5_q0;
  (* dont_touch = "yes" *) reg  cout_V_c_full_n_pass_4_q0;
  always @ (posedge ap_clk) begin
    cout_V_c_full_n_pass_4_q0 <= cout_V_c_full_n_pass_4_out;
  end
  assign cout_V_c_full_n_pass_4_in = cout_V_c_full_n_pass_4_q0;
  (* dont_touch = "yes" *) reg  kernel0_entry12_U0_cout_V_out_write_pass_5_q0;
  always @ (posedge ap_clk) begin
    kernel0_entry12_U0_cout_V_out_write_pass_5_q0 <= kernel0_entry12_U0_cout_V_out_write_pass_5_out;
  end
  assign kernel0_entry12_U0_cout_V_out_write_pass_5_in = kernel0_entry12_U0_cout_V_out_write_pass_5_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper243_U0_fifo_w_out_V_V_din_pass_3_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper243_U0_fifo_w_out_V_V_din_pass_3_q0 <= PE_wrapper243_U0_fifo_w_out_V_V_din_pass_3_out;
  end
  assign PE_wrapper243_U0_fifo_w_out_V_V_din_pass_3_in = PE_wrapper243_U0_fifo_w_out_V_V_din_pass_3_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_7_10_V_V_full_n_pass_2_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_7_10_V_V_full_n_pass_2_q0 <= fifo_w_PE_7_10_V_V_full_n_pass_2_out;
  end
  assign fifo_w_PE_7_10_V_V_full_n_pass_2_in = fifo_w_PE_7_10_V_V_full_n_pass_2_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper243_U0_fifo_w_out_V_V_write_pass_3_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper243_U0_fifo_w_out_V_V_write_pass_3_q0 <= PE_wrapper243_U0_fifo_w_out_V_V_write_pass_3_out;
  end
  assign PE_wrapper243_U0_fifo_w_out_V_V_write_pass_3_in = PE_wrapper243_U0_fifo_w_out_V_V_write_pass_3_q0;
  (* dont_touch = "yes" *) reg [31:0] PE_wrapper243_U0_fifo_cout_drain_out_V_din_pass_3_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper243_U0_fifo_cout_drain_out_V_din_pass_3_q0 <= PE_wrapper243_U0_fifo_cout_drain_out_V_din_pass_3_out;
  end
  assign PE_wrapper243_U0_fifo_cout_drain_out_V_din_pass_3_in = PE_wrapper243_U0_fifo_cout_drain_out_V_din_pass_3_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_PE_7_9_V_full_n_pass_2_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_PE_7_9_V_full_n_pass_2_q0 <= fifo_cout_drain_PE_7_9_V_full_n_pass_2_out;
  end
  assign fifo_cout_drain_PE_7_9_V_full_n_pass_2_in = fifo_cout_drain_PE_7_9_V_full_n_pass_2_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper243_U0_fifo_cout_drain_out_V_write_pass_3_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper243_U0_fifo_cout_drain_out_V_write_pass_3_q0 <= PE_wrapper243_U0_fifo_cout_drain_out_V_write_pass_3_out;
  end
  assign PE_wrapper243_U0_fifo_cout_drain_out_V_write_pass_3_in = PE_wrapper243_U0_fifo_cout_drain_out_V_write_pass_3_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper243_U0_fifo_cin_out_V_V_din_pass_3_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper243_U0_fifo_cin_out_V_V_din_pass_3_q0 <= PE_wrapper243_U0_fifo_cin_out_V_V_din_pass_3_out;
  end
  assign PE_wrapper243_U0_fifo_cin_out_V_V_din_pass_3_in = PE_wrapper243_U0_fifo_cin_out_V_V_din_pass_3_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_8_9_V_V_full_n_pass_2_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_8_9_V_V_full_n_pass_2_q0 <= fifo_cin_PE_8_9_V_V_full_n_pass_2_out;
  end
  assign fifo_cin_PE_8_9_V_V_full_n_pass_2_in = fifo_cin_PE_8_9_V_V_full_n_pass_2_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper243_U0_fifo_cin_out_V_V_write_pass_3_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper243_U0_fifo_cin_out_V_V_write_pass_3_q0 <= PE_wrapper243_U0_fifo_cin_out_V_V_write_pass_3_out;
  end
  assign PE_wrapper243_U0_fifo_cin_out_V_V_write_pass_3_in = PE_wrapper243_U0_fifo_cin_out_V_V_write_pass_3_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper182_U0_fifo_w_out_V_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper182_U0_fifo_w_out_V_V_din_pass_1_q0 <= PE_wrapper182_U0_fifo_w_out_V_V_din_pass_1_out;
  end
  assign PE_wrapper182_U0_fifo_w_out_V_V_din_pass_1_in = PE_wrapper182_U0_fifo_w_out_V_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_2_9_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_2_9_V_V_full_n_pass_0_q0 <= fifo_w_PE_2_9_V_V_full_n_pass_0_out;
  end
  assign fifo_w_PE_2_9_V_V_full_n_pass_0_in = fifo_w_PE_2_9_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper182_U0_fifo_w_out_V_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper182_U0_fifo_w_out_V_V_write_pass_1_q0 <= PE_wrapper182_U0_fifo_w_out_V_V_write_pass_1_out;
  end
  assign PE_wrapper182_U0_fifo_w_out_V_V_write_pass_1_in = PE_wrapper182_U0_fifo_w_out_V_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [63:0] cout_drain_IO_L3_out_U0_fifo_cout_drain_out_V_V_din_pass_2_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L3_out_U0_fifo_cout_drain_out_V_V_din_pass_2_q0 <= cout_drain_IO_L3_out_U0_fifo_cout_drain_out_V_V_din_pass_2_out;
  end
  assign cout_drain_IO_L3_out_U0_fifo_cout_drain_out_V_V_din_pass_2_in = cout_drain_IO_L3_out_U0_fifo_cout_drain_out_V_V_din_pass_2_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_cout_drain_IO_L3_out_serialize_V_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_cout_drain_IO_L3_out_serialize_V_V_full_n_pass_1_q0 <= fifo_cout_drain_cout_drain_IO_L3_out_serialize_V_V_full_n_pass_1_out;
  end
  assign fifo_cout_drain_cout_drain_IO_L3_out_serialize_V_V_full_n_pass_1_in = fifo_cout_drain_cout_drain_IO_L3_out_serialize_V_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg  cout_drain_IO_L3_out_U0_fifo_cout_drain_out_V_V_write_pass_2_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L3_out_U0_fifo_cout_drain_out_V_V_write_pass_2_q0 <= cout_drain_IO_L3_out_U0_fifo_cout_drain_out_V_V_write_pass_2_out;
  end
  assign cout_drain_IO_L3_out_U0_fifo_cout_drain_out_V_V_write_pass_2_in = cout_drain_IO_L3_out_U0_fifo_cout_drain_out_V_V_write_pass_2_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper194_U0_fifo_w_out_V_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper194_U0_fifo_w_out_V_V_din_pass_1_q0 <= PE_wrapper194_U0_fifo_w_out_V_V_din_pass_1_out;
  end
  assign PE_wrapper194_U0_fifo_w_out_V_V_din_pass_1_in = PE_wrapper194_U0_fifo_w_out_V_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_3_9_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_3_9_V_V_full_n_pass_0_q0 <= fifo_w_PE_3_9_V_V_full_n_pass_0_out;
  end
  assign fifo_w_PE_3_9_V_V_full_n_pass_0_in = fifo_w_PE_3_9_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper194_U0_fifo_w_out_V_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper194_U0_fifo_w_out_V_V_write_pass_1_q0 <= PE_wrapper194_U0_fifo_w_out_V_V_write_pass_1_out;
  end
  assign PE_wrapper194_U0_fifo_w_out_V_V_write_pass_1_in = PE_wrapper194_U0_fifo_w_out_V_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper253_U0_fifo_cin_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper253_U0_fifo_cin_out_V_V_din_pass_0_q0 <= PE_wrapper253_U0_fifo_cin_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper253_U0_fifo_cin_out_V_V_din_pass_0_in = PE_wrapper253_U0_fifo_cin_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper253_U0_fifo_cin_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper253_U0_fifo_cin_out_V_V_write_pass_0_q0 <= PE_wrapper253_U0_fifo_cin_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper253_U0_fifo_cin_out_V_V_write_pass_0_in = PE_wrapper253_U0_fifo_cin_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [63:0] cout_drain_IO_L1_out_wrapper471_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper471_U0_fifo_cout_drain_out_V_V_din_pass_0_q0 <= cout_drain_IO_L1_out_wrapper471_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper471_U0_fifo_cout_drain_out_V_V_din_pass_0_in = cout_drain_IO_L1_out_wrapper471_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  cout_drain_IO_L1_out_wrapper471_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper471_U0_fifo_cout_drain_out_V_V_write_pass_0_q0 <= cout_drain_IO_L1_out_wrapper471_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper471_U0_fifo_cout_drain_out_V_V_write_pass_0_in = cout_drain_IO_L1_out_wrapper471_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_PE_5_8_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_PE_5_8_V_full_n_pass_0_q0 <= fifo_cout_drain_PE_5_8_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_PE_5_8_V_full_n_pass_0_in = fifo_cout_drain_PE_5_8_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper242_U0_fifo_w_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper242_U0_fifo_w_out_V_V_din_pass_0_q0 <= PE_wrapper242_U0_fifo_w_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper242_U0_fifo_w_out_V_V_din_pass_0_in = PE_wrapper242_U0_fifo_w_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper242_U0_fifo_w_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper242_U0_fifo_w_out_V_V_write_pass_0_q0 <= PE_wrapper242_U0_fifo_w_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper242_U0_fifo_w_out_V_V_write_pass_0_in = PE_wrapper242_U0_fifo_w_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper230_U0_fifo_w_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper230_U0_fifo_w_out_V_V_din_pass_0_q0 <= PE_wrapper230_U0_fifo_w_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper230_U0_fifo_w_out_V_V_din_pass_0_in = PE_wrapper230_U0_fifo_w_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper230_U0_fifo_w_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper230_U0_fifo_w_out_V_V_write_pass_0_q0 <= PE_wrapper230_U0_fifo_w_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper230_U0_fifo_w_out_V_V_write_pass_0_in = PE_wrapper230_U0_fifo_w_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [63:0] cout_drain_IO_L1_out_wrapper506_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper506_U0_fifo_cout_drain_out_V_V_din_pass_0_q0 <= cout_drain_IO_L1_out_wrapper506_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper506_U0_fifo_cout_drain_out_V_V_din_pass_0_in = cout_drain_IO_L1_out_wrapper506_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  cout_drain_IO_L1_out_wrapper506_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper506_U0_fifo_cout_drain_out_V_V_write_pass_0_q0 <= cout_drain_IO_L1_out_wrapper506_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper506_U0_fifo_cout_drain_out_V_V_write_pass_0_in = cout_drain_IO_L1_out_wrapper506_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper252_U0_fifo_cin_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper252_U0_fifo_cin_out_V_V_din_pass_0_q0 <= PE_wrapper252_U0_fifo_cin_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper252_U0_fifo_cin_out_V_V_din_pass_0_in = PE_wrapper252_U0_fifo_cin_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper252_U0_fifo_cin_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper252_U0_fifo_cin_out_V_V_write_pass_0_q0 <= PE_wrapper252_U0_fifo_cin_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper252_U0_fifo_cin_out_V_V_write_pass_0_in = PE_wrapper252_U0_fifo_cin_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_7_6_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_7_6_V_V_full_n_pass_0_q0 <= fifo_cin_PE_7_6_V_V_full_n_pass_0_out;
  end
  assign fifo_cin_PE_7_6_V_V_full_n_pass_0_in = fifo_cin_PE_7_6_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper254_U0_fifo_w_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper254_U0_fifo_w_out_V_V_din_pass_0_q0 <= PE_wrapper254_U0_fifo_w_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper254_U0_fifo_w_out_V_V_din_pass_0_in = PE_wrapper254_U0_fifo_w_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper254_U0_fifo_w_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper254_U0_fifo_w_out_V_V_write_pass_0_q0 <= PE_wrapper254_U0_fifo_w_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper254_U0_fifo_w_out_V_V_write_pass_0_in = PE_wrapper254_U0_fifo_w_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_cout_drain_IO_L1_out_8_9_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_cout_drain_IO_L1_out_8_9_V_V_full_n_pass_0_q0 <= fifo_cout_drain_cout_drain_IO_L1_out_8_9_V_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_cout_drain_IO_L1_out_8_9_V_V_full_n_pass_0_in = fifo_cout_drain_cout_drain_IO_L1_out_8_9_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_6_8_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_6_8_V_V_full_n_pass_0_q0 <= fifo_w_PE_6_8_V_V_full_n_pass_0_out;
  end
  assign fifo_w_PE_6_8_V_V_full_n_pass_0_in = fifo_w_PE_6_8_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_7_7_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_7_7_V_V_full_n_pass_0_q0 <= fifo_cin_PE_7_7_V_V_full_n_pass_0_out;
  end
  assign fifo_cin_PE_7_7_V_V_full_n_pass_0_in = fifo_cin_PE_7_7_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_8_6_V_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_8_6_V_V_full_n_pass_1_q0 <= fifo_w_PE_8_6_V_V_full_n_pass_1_out;
  end
  assign fifo_w_PE_8_6_V_V_full_n_pass_1_in = fifo_w_PE_8_6_V_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_cout_drain_IO_L1_out_7_9_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_cout_drain_IO_L1_out_7_9_V_V_full_n_pass_0_q0 <= fifo_cout_drain_cout_drain_IO_L1_out_7_9_V_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_cout_drain_IO_L1_out_7_9_V_V_full_n_pass_0_in = fifo_cout_drain_cout_drain_IO_L1_out_7_9_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg [63:0] cout_drain_IO_L1_out_wrapper487_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper487_U0_fifo_cout_drain_out_V_V_din_pass_0_q0 <= cout_drain_IO_L1_out_wrapper487_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper487_U0_fifo_cout_drain_out_V_V_din_pass_0_in = cout_drain_IO_L1_out_wrapper487_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  cout_drain_IO_L1_out_wrapper487_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper487_U0_fifo_cout_drain_out_V_V_write_pass_0_q0 <= cout_drain_IO_L1_out_wrapper487_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper487_U0_fifo_cout_drain_out_V_V_write_pass_0_in = cout_drain_IO_L1_out_wrapper487_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_PE_4_8_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_PE_4_8_V_full_n_pass_0_q0 <= fifo_cout_drain_PE_4_8_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_PE_4_8_V_full_n_pass_0_in = fifo_cout_drain_PE_4_8_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_6_8_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_6_8_V_V_full_n_pass_0_q0 <= fifo_cin_PE_6_8_V_V_full_n_pass_0_out;
  end
  assign fifo_cin_PE_6_8_V_V_full_n_pass_0_in = fifo_cin_PE_6_8_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_7_6_V_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_7_6_V_V_full_n_pass_1_q0 <= fifo_w_PE_7_6_V_V_full_n_pass_1_out;
  end
  assign fifo_w_PE_7_6_V_V_full_n_pass_1_in = fifo_w_PE_7_6_V_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper254_U0_fifo_cin_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper254_U0_fifo_cin_out_V_V_din_pass_0_q0 <= PE_wrapper254_U0_fifo_cin_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper254_U0_fifo_cin_out_V_V_din_pass_0_in = PE_wrapper254_U0_fifo_cin_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper254_U0_fifo_cin_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper254_U0_fifo_cin_out_V_V_write_pass_0_q0 <= PE_wrapper254_U0_fifo_cin_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper254_U0_fifo_cin_out_V_V_write_pass_0_in = PE_wrapper254_U0_fifo_cin_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_cout_drain_IO_L1_out_6_9_V_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_cout_drain_IO_L1_out_6_9_V_V_full_n_pass_1_q0 <= fifo_cout_drain_cout_drain_IO_L1_out_6_9_V_V_full_n_pass_1_out;
  end
  assign fifo_cout_drain_cout_drain_IO_L1_out_6_9_V_V_full_n_pass_1_in = fifo_cout_drain_cout_drain_IO_L1_out_6_9_V_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg  ap_done_Boundary_X4Y10_To_X6Y10_q0;
  always @ (posedge ap_clk) begin
    ap_done_Boundary_X4Y10_To_X6Y10_q0 <= ap_done_Boundary_X4Y10_To_X6Y10_out;
  end
  assign ap_done_Boundary_X4Y10_To_X6Y10_in = ap_done_Boundary_X4Y10_To_X6Y10_q0;
  (* dont_touch = "yes" *) reg  ap_start_Boundary_X4Y12_To_X6Y12_q0;
  always @ (posedge ap_clk) begin
    ap_start_Boundary_X4Y12_To_X6Y12_q0 <= ap_start_Boundary_X4Y12_To_X6Y12_out;
  end
  assign ap_start_Boundary_X4Y12_To_X6Y12_in = ap_start_Boundary_X4Y12_To_X6Y12_q0;
  (* dont_touch = "yes" *) reg  ap_rst_n_Boundary_X4Y12_To_X6Y12_q0;
  always @ (posedge ap_clk) begin
    ap_rst_n_Boundary_X4Y12_To_X6Y12_q0 <= ap_rst_n_Boundary_X4Y12_To_X6Y12_out;
  end
  assign ap_rst_n_Boundary_X4Y12_To_X6Y12_in = ap_rst_n_Boundary_X4Y12_To_X6Y12_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper242_U0_fifo_w_out_V_V_din_pass_2_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper242_U0_fifo_w_out_V_V_din_pass_2_q0 <= PE_wrapper242_U0_fifo_w_out_V_V_din_pass_2_out;
  end
  assign PE_wrapper242_U0_fifo_w_out_V_V_din_pass_2_in = PE_wrapper242_U0_fifo_w_out_V_V_din_pass_2_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_7_9_V_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_7_9_V_V_full_n_pass_1_q0 <= fifo_w_PE_7_9_V_V_full_n_pass_1_out;
  end
  assign fifo_w_PE_7_9_V_V_full_n_pass_1_in = fifo_w_PE_7_9_V_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper242_U0_fifo_w_out_V_V_write_pass_2_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper242_U0_fifo_w_out_V_V_write_pass_2_q0 <= PE_wrapper242_U0_fifo_w_out_V_V_write_pass_2_out;
  end
  assign PE_wrapper242_U0_fifo_w_out_V_V_write_pass_2_in = PE_wrapper242_U0_fifo_w_out_V_V_write_pass_2_q0;
  (* dont_touch = "yes" *) reg [63:0] cout_drain_IO_L1_out_wrapper474_U0_fifo_cout_drain_out_V_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper474_U0_fifo_cout_drain_out_V_V_din_pass_1_q0 <= cout_drain_IO_L1_out_wrapper474_U0_fifo_cout_drain_out_V_V_din_pass_1_out;
  end
  assign cout_drain_IO_L1_out_wrapper474_U0_fifo_cout_drain_out_V_V_din_pass_1_in = cout_drain_IO_L1_out_wrapper474_U0_fifo_cout_drain_out_V_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_cout_drain_IO_L1_out_6_4_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_cout_drain_IO_L1_out_6_4_V_V_full_n_pass_0_q0 <= fifo_cout_drain_cout_drain_IO_L1_out_6_4_V_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_cout_drain_IO_L1_out_6_4_V_V_full_n_pass_0_in = fifo_cout_drain_cout_drain_IO_L1_out_6_4_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  cout_drain_IO_L1_out_wrapper474_U0_fifo_cout_drain_out_V_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper474_U0_fifo_cout_drain_out_V_V_write_pass_1_q0 <= cout_drain_IO_L1_out_wrapper474_U0_fifo_cout_drain_out_V_V_write_pass_1_out;
  end
  assign cout_drain_IO_L1_out_wrapper474_U0_fifo_cout_drain_out_V_V_write_pass_1_in = cout_drain_IO_L1_out_wrapper474_U0_fifo_cout_drain_out_V_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [63:0] cout_drain_IO_L1_out_wrapper458_U0_fifo_cout_drain_out_V_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper458_U0_fifo_cout_drain_out_V_V_din_pass_1_q0 <= cout_drain_IO_L1_out_wrapper458_U0_fifo_cout_drain_out_V_V_din_pass_1_out;
  end
  assign cout_drain_IO_L1_out_wrapper458_U0_fifo_cout_drain_out_V_V_din_pass_1_in = cout_drain_IO_L1_out_wrapper458_U0_fifo_cout_drain_out_V_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_cout_drain_IO_L1_out_5_4_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_cout_drain_IO_L1_out_5_4_V_V_full_n_pass_0_q0 <= fifo_cout_drain_cout_drain_IO_L1_out_5_4_V_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_cout_drain_IO_L1_out_5_4_V_V_full_n_pass_0_in = fifo_cout_drain_cout_drain_IO_L1_out_5_4_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  cout_drain_IO_L1_out_wrapper458_U0_fifo_cout_drain_out_V_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper458_U0_fifo_cout_drain_out_V_V_write_pass_1_q0 <= cout_drain_IO_L1_out_wrapper458_U0_fifo_cout_drain_out_V_V_write_pass_1_out;
  end
  assign cout_drain_IO_L1_out_wrapper458_U0_fifo_cout_drain_out_V_V_write_pass_1_in = cout_drain_IO_L1_out_wrapper458_U0_fifo_cout_drain_out_V_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper231_U0_fifo_cin_out_V_V_din_pass_4_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper231_U0_fifo_cin_out_V_V_din_pass_4_q0 <= PE_wrapper231_U0_fifo_cin_out_V_V_din_pass_4_out;
  end
  assign PE_wrapper231_U0_fifo_cin_out_V_V_din_pass_4_in = PE_wrapper231_U0_fifo_cin_out_V_V_din_pass_4_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_7_9_V_V_full_n_pass_3_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_7_9_V_V_full_n_pass_3_q0 <= fifo_cin_PE_7_9_V_V_full_n_pass_3_out;
  end
  assign fifo_cin_PE_7_9_V_V_full_n_pass_3_in = fifo_cin_PE_7_9_V_V_full_n_pass_3_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper231_U0_fifo_cin_out_V_V_write_pass_4_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper231_U0_fifo_cin_out_V_V_write_pass_4_q0 <= PE_wrapper231_U0_fifo_cin_out_V_V_write_pass_4_out;
  end
  assign PE_wrapper231_U0_fifo_cin_out_V_V_write_pass_4_in = PE_wrapper231_U0_fifo_cin_out_V_V_write_pass_4_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper217_U0_fifo_w_out_V_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper217_U0_fifo_w_out_V_V_din_pass_1_q0 <= PE_wrapper217_U0_fifo_w_out_V_V_din_pass_1_out;
  end
  assign PE_wrapper217_U0_fifo_w_out_V_V_din_pass_1_in = PE_wrapper217_U0_fifo_w_out_V_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_5_8_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_5_8_V_V_full_n_pass_0_q0 <= fifo_w_PE_5_8_V_V_full_n_pass_0_out;
  end
  assign fifo_w_PE_5_8_V_V_full_n_pass_0_in = fifo_w_PE_5_8_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper217_U0_fifo_w_out_V_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper217_U0_fifo_w_out_V_V_write_pass_1_q0 <= PE_wrapper217_U0_fifo_w_out_V_V_write_pass_1_out;
  end
  assign PE_wrapper217_U0_fifo_w_out_V_V_write_pass_1_in = PE_wrapper217_U0_fifo_w_out_V_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_1_7_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_1_7_V_V_full_n_pass_0_q0 <= fifo_w_PE_1_7_V_V_full_n_pass_0_out;
  end
  assign fifo_w_PE_1_7_V_V_full_n_pass_0_in = fifo_w_PE_1_7_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper193_U0_fifo_w_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper193_U0_fifo_w_out_V_V_din_pass_0_q0 <= PE_wrapper193_U0_fifo_w_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper193_U0_fifo_w_out_V_V_din_pass_0_in = PE_wrapper193_U0_fifo_w_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper193_U0_fifo_w_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper193_U0_fifo_w_out_V_V_write_pass_0_q0 <= PE_wrapper193_U0_fifo_w_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper193_U0_fifo_w_out_V_V_write_pass_0_in = PE_wrapper193_U0_fifo_w_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper181_U0_fifo_w_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper181_U0_fifo_w_out_V_V_din_pass_0_q0 <= PE_wrapper181_U0_fifo_w_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper181_U0_fifo_w_out_V_V_din_pass_0_in = PE_wrapper181_U0_fifo_w_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper181_U0_fifo_w_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper181_U0_fifo_w_out_V_V_write_pass_0_q0 <= PE_wrapper181_U0_fifo_w_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper181_U0_fifo_w_out_V_V_write_pass_0_in = PE_wrapper181_U0_fifo_w_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [63:0] cout_drain_IO_L2_out561_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L2_out561_U0_fifo_cout_drain_out_V_V_din_pass_0_q0 <= cout_drain_IO_L2_out561_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  end
  assign cout_drain_IO_L2_out561_U0_fifo_cout_drain_out_V_V_din_pass_0_in = cout_drain_IO_L2_out561_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  cout_drain_IO_L2_out561_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L2_out561_U0_fifo_cout_drain_out_V_V_write_pass_0_q0 <= cout_drain_IO_L2_out561_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  end
  assign cout_drain_IO_L2_out561_U0_fifo_cout_drain_out_V_V_write_pass_0_in = cout_drain_IO_L2_out561_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper169_U0_fifo_w_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper169_U0_fifo_w_out_V_V_din_pass_0_q0 <= PE_wrapper169_U0_fifo_w_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper169_U0_fifo_w_out_V_V_din_pass_0_in = PE_wrapper169_U0_fifo_w_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper169_U0_fifo_w_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper169_U0_fifo_w_out_V_V_write_pass_0_q0 <= PE_wrapper169_U0_fifo_w_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper169_U0_fifo_w_out_V_V_write_pass_0_in = PE_wrapper169_U0_fifo_w_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_cin_IO_L2_in_7_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_cin_IO_L2_in_7_V_V_full_n_pass_0_q0 <= fifo_cin_cin_IO_L2_in_7_V_V_full_n_pass_0_out;
  end
  assign fifo_cin_cin_IO_L2_in_7_V_V_full_n_pass_0_in = fifo_cin_cin_IO_L2_in_7_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper205_U0_fifo_cin_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper205_U0_fifo_cin_out_V_V_din_pass_0_q0 <= PE_wrapper205_U0_fifo_cin_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper205_U0_fifo_cin_out_V_V_din_pass_0_in = PE_wrapper205_U0_fifo_cin_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper205_U0_fifo_cin_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper205_U0_fifo_cin_out_V_V_write_pass_0_q0 <= PE_wrapper205_U0_fifo_cin_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper205_U0_fifo_cin_out_V_V_write_pass_0_in = PE_wrapper205_U0_fifo_cin_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_cout_drain_IO_L1_out_7_4_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_cout_drain_IO_L1_out_7_4_V_V_full_n_pass_0_q0 <= fifo_cout_drain_cout_drain_IO_L1_out_7_4_V_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_cout_drain_IO_L1_out_7_4_V_V_full_n_pass_0_in = fifo_cout_drain_cout_drain_IO_L1_out_7_4_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] cin_IO_L2_in131_U0_fifo_cin_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    cin_IO_L2_in131_U0_fifo_cin_out_V_V_din_pass_0_q0 <= cin_IO_L2_in131_U0_fifo_cin_out_V_V_din_pass_0_out;
  end
  assign cin_IO_L2_in131_U0_fifo_cin_out_V_V_din_pass_0_in = cin_IO_L2_in131_U0_fifo_cin_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  cin_IO_L2_in131_U0_fifo_cin_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    cin_IO_L2_in131_U0_fifo_cin_out_V_V_write_pass_0_q0 <= cin_IO_L2_in131_U0_fifo_cin_out_V_V_write_pass_0_out;
  end
  assign cin_IO_L2_in131_U0_fifo_cin_out_V_V_write_pass_0_in = cin_IO_L2_in131_U0_fifo_cin_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_0_7_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_0_7_V_V_full_n_pass_0_q0 <= fifo_w_PE_0_7_V_V_full_n_pass_0_out;
  end
  assign fifo_w_PE_0_7_V_V_full_n_pass_0_in = fifo_w_PE_0_7_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper157_U0_fifo_w_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper157_U0_fifo_w_out_V_V_din_pass_0_q0 <= PE_wrapper157_U0_fifo_w_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper157_U0_fifo_w_out_V_V_din_pass_0_in = PE_wrapper157_U0_fifo_w_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper157_U0_fifo_w_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper157_U0_fifo_w_out_V_V_write_pass_0_q0 <= PE_wrapper157_U0_fifo_w_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper157_U0_fifo_w_out_V_V_write_pass_0_in = PE_wrapper157_U0_fifo_w_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_3_7_V_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_3_7_V_V_full_n_pass_1_q0 <= fifo_w_PE_3_7_V_V_full_n_pass_1_out;
  end
  assign fifo_w_PE_3_7_V_V_full_n_pass_1_in = fifo_w_PE_3_7_V_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_cout_drain_IO_L2_out_8_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_cout_drain_IO_L2_out_8_V_V_full_n_pass_0_q0 <= fifo_cout_drain_cout_drain_IO_L2_out_8_V_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_cout_drain_IO_L2_out_8_V_V_full_n_pass_0_in = fifo_cout_drain_cout_drain_IO_L2_out_8_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg [63:0] cout_drain_IO_L3_out_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L3_out_U0_fifo_cout_drain_out_V_V_din_pass_0_q0 <= cout_drain_IO_L3_out_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  end
  assign cout_drain_IO_L3_out_U0_fifo_cout_drain_out_V_V_din_pass_0_in = cout_drain_IO_L3_out_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  cout_drain_IO_L3_out_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L3_out_U0_fifo_cout_drain_out_V_V_write_pass_0_q0 <= cout_drain_IO_L3_out_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  end
  assign cout_drain_IO_L3_out_U0_fifo_cout_drain_out_V_V_write_pass_0_in = cout_drain_IO_L3_out_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_2_7_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_2_7_V_V_full_n_pass_0_q0 <= fifo_w_PE_2_7_V_V_full_n_pass_0_out;
  end
  assign fifo_w_PE_2_7_V_V_full_n_pass_0_in = fifo_w_PE_2_7_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg [31:0] PE_wrapper205_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper205_U0_fifo_cout_drain_out_V_din_pass_0_q0 <= PE_wrapper205_U0_fifo_cout_drain_out_V_din_pass_0_out;
  end
  assign PE_wrapper205_U0_fifo_cout_drain_out_V_din_pass_0_in = PE_wrapper205_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper205_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper205_U0_fifo_cout_drain_out_V_write_pass_0_q0 <= PE_wrapper205_U0_fifo_cout_drain_out_V_write_pass_0_out;
  end
  assign PE_wrapper205_U0_fifo_cout_drain_out_V_write_pass_0_in = PE_wrapper205_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper205_U0_fifo_w_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper205_U0_fifo_w_out_V_V_din_pass_0_q0 <= PE_wrapper205_U0_fifo_w_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper205_U0_fifo_w_out_V_V_din_pass_0_in = PE_wrapper205_U0_fifo_w_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper205_U0_fifo_w_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper205_U0_fifo_w_out_V_V_write_pass_0_q0 <= PE_wrapper205_U0_fifo_w_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper205_U0_fifo_w_out_V_V_write_pass_0_in = PE_wrapper205_U0_fifo_w_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_4_7_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_4_7_V_V_full_n_pass_0_q0 <= fifo_w_PE_4_7_V_V_full_n_pass_0_out;
  end
  assign fifo_w_PE_4_7_V_V_full_n_pass_0_in = fifo_w_PE_4_7_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_cout_drain_IO_L2_out_0_V_V_full_n_pass_3_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_cout_drain_IO_L2_out_0_V_V_full_n_pass_3_q0 <= fifo_cout_drain_cout_drain_IO_L2_out_0_V_V_full_n_pass_3_out;
  end
  assign fifo_cout_drain_cout_drain_IO_L2_out_0_V_V_full_n_pass_3_in = fifo_cout_drain_cout_drain_IO_L2_out_0_V_V_full_n_pass_3_q0;
  (* dont_touch = "yes" *) reg  ap_done_Boundary_X6Y8_To_X8Y8_q0;
  always @ (posedge ap_clk) begin
    ap_done_Boundary_X6Y8_To_X8Y8_q0 <= ap_done_Boundary_X6Y8_To_X8Y8_out;
  end
  assign ap_done_Boundary_X6Y8_To_X8Y8_in = ap_done_Boundary_X6Y8_To_X8Y8_q0;
  (* dont_touch = "yes" *) reg  ap_start_Boundary_X6Y10_To_X8Y10_q0;
  always @ (posedge ap_clk) begin
    ap_start_Boundary_X6Y10_To_X8Y10_q0 <= ap_start_Boundary_X6Y10_To_X8Y10_out;
  end
  assign ap_start_Boundary_X6Y10_To_X8Y10_in = ap_start_Boundary_X6Y10_To_X8Y10_q0;
  (* dont_touch = "yes" *) reg  ap_rst_n_Boundary_X6Y10_To_X8Y10_q0;
  always @ (posedge ap_clk) begin
    ap_rst_n_Boundary_X6Y10_To_X8Y10_q0 <= ap_rst_n_Boundary_X6Y10_To_X8Y10_out;
  end
  assign ap_rst_n_Boundary_X6Y10_To_X8Y10_in = ap_rst_n_Boundary_X6Y10_To_X8Y10_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper242_U0_fifo_w_out_V_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper242_U0_fifo_w_out_V_V_din_pass_1_q0 <= PE_wrapper242_U0_fifo_w_out_V_V_din_pass_1_out;
  end
  assign PE_wrapper242_U0_fifo_w_out_V_V_din_pass_1_in = PE_wrapper242_U0_fifo_w_out_V_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_7_9_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_7_9_V_V_full_n_pass_0_q0 <= fifo_w_PE_7_9_V_V_full_n_pass_0_out;
  end
  assign fifo_w_PE_7_9_V_V_full_n_pass_0_in = fifo_w_PE_7_9_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper242_U0_fifo_w_out_V_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper242_U0_fifo_w_out_V_V_write_pass_1_q0 <= PE_wrapper242_U0_fifo_w_out_V_V_write_pass_1_out;
  end
  assign PE_wrapper242_U0_fifo_w_out_V_V_write_pass_1_in = PE_wrapper242_U0_fifo_w_out_V_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper231_U0_fifo_cin_out_V_V_din_pass_3_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper231_U0_fifo_cin_out_V_V_din_pass_3_q0 <= PE_wrapper231_U0_fifo_cin_out_V_V_din_pass_3_out;
  end
  assign PE_wrapper231_U0_fifo_cin_out_V_V_din_pass_3_in = PE_wrapper231_U0_fifo_cin_out_V_V_din_pass_3_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_7_9_V_V_full_n_pass_2_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_7_9_V_V_full_n_pass_2_q0 <= fifo_cin_PE_7_9_V_V_full_n_pass_2_out;
  end
  assign fifo_cin_PE_7_9_V_V_full_n_pass_2_in = fifo_cin_PE_7_9_V_V_full_n_pass_2_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper231_U0_fifo_cin_out_V_V_write_pass_3_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper231_U0_fifo_cin_out_V_V_write_pass_3_q0 <= PE_wrapper231_U0_fifo_cin_out_V_V_write_pass_3_out;
  end
  assign PE_wrapper231_U0_fifo_cin_out_V_V_write_pass_3_in = PE_wrapper231_U0_fifo_cin_out_V_V_write_pass_3_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper158_U0_fifo_w_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper158_U0_fifo_w_out_V_V_din_pass_0_q0 <= PE_wrapper158_U0_fifo_w_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper158_U0_fifo_w_out_V_V_din_pass_0_in = PE_wrapper158_U0_fifo_w_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper158_U0_fifo_w_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper158_U0_fifo_w_out_V_V_write_pass_0_q0 <= PE_wrapper158_U0_fifo_w_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper158_U0_fifo_w_out_V_V_write_pass_0_in = PE_wrapper158_U0_fifo_w_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_3_8_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_3_8_V_V_full_n_pass_0_q0 <= fifo_w_PE_3_8_V_V_full_n_pass_0_out;
  end
  assign fifo_w_PE_3_8_V_V_full_n_pass_0_in = fifo_w_PE_3_8_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper170_U0_fifo_w_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper170_U0_fifo_w_out_V_V_din_pass_0_q0 <= PE_wrapper170_U0_fifo_w_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper170_U0_fifo_w_out_V_V_din_pass_0_in = PE_wrapper170_U0_fifo_w_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper170_U0_fifo_w_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper170_U0_fifo_w_out_V_V_write_pass_0_q0 <= PE_wrapper170_U0_fifo_w_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper170_U0_fifo_w_out_V_V_write_pass_0_in = PE_wrapper170_U0_fifo_w_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_cout_drain_IO_L2_out_9_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_cout_drain_IO_L2_out_9_V_V_full_n_pass_0_q0 <= fifo_cout_drain_cout_drain_IO_L2_out_9_V_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_cout_drain_IO_L2_out_9_V_V_full_n_pass_0_in = fifo_cout_drain_cout_drain_IO_L2_out_9_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_2_8_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_2_8_V_V_full_n_pass_0_q0 <= fifo_w_PE_2_8_V_V_full_n_pass_0_out;
  end
  assign fifo_w_PE_2_8_V_V_full_n_pass_0_in = fifo_w_PE_2_8_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper206_U0_fifo_w_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper206_U0_fifo_w_out_V_V_din_pass_0_q0 <= PE_wrapper206_U0_fifo_w_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper206_U0_fifo_w_out_V_V_din_pass_0_in = PE_wrapper206_U0_fifo_w_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper206_U0_fifo_w_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper206_U0_fifo_w_out_V_V_write_pass_0_q0 <= PE_wrapper206_U0_fifo_w_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper206_U0_fifo_w_out_V_V_write_pass_0_in = PE_wrapper206_U0_fifo_w_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] cin_IO_L2_in132_U0_fifo_cin_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    cin_IO_L2_in132_U0_fifo_cin_out_V_V_din_pass_0_q0 <= cin_IO_L2_in132_U0_fifo_cin_out_V_V_din_pass_0_out;
  end
  assign cin_IO_L2_in132_U0_fifo_cin_out_V_V_din_pass_0_in = cin_IO_L2_in132_U0_fifo_cin_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  cin_IO_L2_in132_U0_fifo_cin_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    cin_IO_L2_in132_U0_fifo_cin_out_V_V_write_pass_0_q0 <= cin_IO_L2_in132_U0_fifo_cin_out_V_V_write_pass_0_out;
  end
  assign cin_IO_L2_in132_U0_fifo_cin_out_V_V_write_pass_0_in = cin_IO_L2_in132_U0_fifo_cin_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [31:0] PE_wrapper218_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper218_U0_fifo_cout_drain_out_V_din_pass_0_q0 <= PE_wrapper218_U0_fifo_cout_drain_out_V_din_pass_0_out;
  end
  assign PE_wrapper218_U0_fifo_cout_drain_out_V_din_pass_0_in = PE_wrapper218_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper218_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper218_U0_fifo_cout_drain_out_V_write_pass_0_q0 <= PE_wrapper218_U0_fifo_cout_drain_out_V_write_pass_0_out;
  end
  assign PE_wrapper218_U0_fifo_cout_drain_out_V_write_pass_0_in = PE_wrapper218_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_cout_drain_IO_L1_out_8_4_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_cout_drain_IO_L1_out_8_4_V_V_full_n_pass_0_q0 <= fifo_cout_drain_cout_drain_IO_L1_out_8_4_V_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_cout_drain_IO_L1_out_8_4_V_V_full_n_pass_0_in = fifo_cout_drain_cout_drain_IO_L1_out_8_4_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_1_8_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_1_8_V_V_full_n_pass_0_q0 <= fifo_w_PE_1_8_V_V_full_n_pass_0_out;
  end
  assign fifo_w_PE_1_8_V_V_full_n_pass_0_in = fifo_w_PE_1_8_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_5_8_V_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_5_8_V_V_full_n_pass_1_q0 <= fifo_w_PE_5_8_V_V_full_n_pass_1_out;
  end
  assign fifo_w_PE_5_8_V_V_full_n_pass_1_in = fifo_w_PE_5_8_V_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_cin_IO_L2_in_8_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_cin_IO_L2_in_8_V_V_full_n_pass_0_q0 <= fifo_cin_cin_IO_L2_in_8_V_V_full_n_pass_0_out;
  end
  assign fifo_cin_cin_IO_L2_in_8_V_V_full_n_pass_0_in = fifo_cin_cin_IO_L2_in_8_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_0_8_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_0_8_V_V_full_n_pass_0_q0 <= fifo_w_PE_0_8_V_V_full_n_pass_0_out;
  end
  assign fifo_w_PE_0_8_V_V_full_n_pass_0_in = fifo_w_PE_0_8_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper182_U0_fifo_w_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper182_U0_fifo_w_out_V_V_din_pass_0_q0 <= PE_wrapper182_U0_fifo_w_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper182_U0_fifo_w_out_V_V_din_pass_0_in = PE_wrapper182_U0_fifo_w_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper182_U0_fifo_w_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper182_U0_fifo_w_out_V_V_write_pass_0_q0 <= PE_wrapper182_U0_fifo_w_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper182_U0_fifo_w_out_V_V_write_pass_0_in = PE_wrapper182_U0_fifo_w_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [63:0] cout_drain_IO_L2_out560_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L2_out560_U0_fifo_cout_drain_out_V_V_din_pass_0_q0 <= cout_drain_IO_L2_out560_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  end
  assign cout_drain_IO_L2_out560_U0_fifo_cout_drain_out_V_V_din_pass_0_in = cout_drain_IO_L2_out560_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  cout_drain_IO_L2_out560_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L2_out560_U0_fifo_cout_drain_out_V_V_write_pass_0_q0 <= cout_drain_IO_L2_out560_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  end
  assign cout_drain_IO_L2_out560_U0_fifo_cout_drain_out_V_V_write_pass_0_in = cout_drain_IO_L2_out560_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_4_8_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_4_8_V_V_full_n_pass_0_q0 <= fifo_w_PE_4_8_V_V_full_n_pass_0_out;
  end
  assign fifo_w_PE_4_8_V_V_full_n_pass_0_in = fifo_w_PE_4_8_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper218_U0_fifo_w_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper218_U0_fifo_w_out_V_V_din_pass_0_q0 <= PE_wrapper218_U0_fifo_w_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper218_U0_fifo_w_out_V_V_din_pass_0_in = PE_wrapper218_U0_fifo_w_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper218_U0_fifo_w_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper218_U0_fifo_w_out_V_V_write_pass_0_q0 <= PE_wrapper218_U0_fifo_w_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper218_U0_fifo_w_out_V_V_write_pass_0_in = PE_wrapper218_U0_fifo_w_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [31:0] PE_wrapper206_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper206_U0_fifo_cout_drain_out_V_din_pass_0_q0 <= PE_wrapper206_U0_fifo_cout_drain_out_V_din_pass_0_out;
  end
  assign PE_wrapper206_U0_fifo_cout_drain_out_V_din_pass_0_in = PE_wrapper206_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper206_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper206_U0_fifo_cout_drain_out_V_write_pass_0_q0 <= PE_wrapper206_U0_fifo_cout_drain_out_V_write_pass_0_out;
  end
  assign PE_wrapper206_U0_fifo_cout_drain_out_V_write_pass_0_in = PE_wrapper206_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper218_U0_fifo_cin_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper218_U0_fifo_cin_out_V_V_din_pass_0_q0 <= PE_wrapper218_U0_fifo_cin_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper218_U0_fifo_cin_out_V_V_din_pass_0_in = PE_wrapper218_U0_fifo_cin_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper218_U0_fifo_cin_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper218_U0_fifo_cin_out_V_V_write_pass_0_q0 <= PE_wrapper218_U0_fifo_cin_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper218_U0_fifo_cin_out_V_V_write_pass_0_in = PE_wrapper218_U0_fifo_cin_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper194_U0_fifo_w_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper194_U0_fifo_w_out_V_V_din_pass_0_q0 <= PE_wrapper194_U0_fifo_w_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper194_U0_fifo_w_out_V_V_din_pass_0_in = PE_wrapper194_U0_fifo_w_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper194_U0_fifo_w_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper194_U0_fifo_w_out_V_V_write_pass_0_q0 <= PE_wrapper194_U0_fifo_w_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper194_U0_fifo_w_out_V_V_write_pass_0_in = PE_wrapper194_U0_fifo_w_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  ap_done_Boundary_X6Y10_To_X8Y10_q0;
  always @ (posedge ap_clk) begin
    ap_done_Boundary_X6Y10_To_X8Y10_q0 <= ap_done_Boundary_X6Y10_To_X8Y10_out;
  end
  assign ap_done_Boundary_X6Y10_To_X8Y10_in = ap_done_Boundary_X6Y10_To_X8Y10_q0;
  (* dont_touch = "yes" *) reg  ap_start_Boundary_X6Y12_To_X8Y12_q0;
  always @ (posedge ap_clk) begin
    ap_start_Boundary_X6Y12_To_X8Y12_q0 <= ap_start_Boundary_X6Y12_To_X8Y12_out;
  end
  assign ap_start_Boundary_X6Y12_To_X8Y12_in = ap_start_Boundary_X6Y12_To_X8Y12_q0;
  (* dont_touch = "yes" *) reg  ap_rst_n_Boundary_X6Y12_To_X8Y12_q0;
  always @ (posedge ap_clk) begin
    ap_rst_n_Boundary_X6Y12_To_X8Y12_q0 <= ap_rst_n_Boundary_X6Y12_To_X8Y12_out;
  end
  assign ap_rst_n_Boundary_X6Y12_To_X8Y12_in = ap_rst_n_Boundary_X6Y12_To_X8Y12_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper256_U0_fifo_cin_out_V_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper256_U0_fifo_cin_out_V_V_din_pass_1_q0 <= PE_wrapper256_U0_fifo_cin_out_V_V_din_pass_1_out;
  end
  assign PE_wrapper256_U0_fifo_cin_out_V_V_din_pass_1_in = PE_wrapper256_U0_fifo_cin_out_V_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_9_10_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_9_10_V_V_full_n_pass_0_q0 <= fifo_cin_PE_9_10_V_V_full_n_pass_0_out;
  end
  assign fifo_cin_PE_9_10_V_V_full_n_pass_0_in = fifo_cin_PE_9_10_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper256_U0_fifo_cin_out_V_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper256_U0_fifo_cin_out_V_V_write_pass_1_q0 <= PE_wrapper256_U0_fifo_cin_out_V_V_write_pass_1_out;
  end
  assign PE_wrapper256_U0_fifo_cin_out_V_V_write_pass_1_in = PE_wrapper256_U0_fifo_cin_out_V_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper257_U0_fifo_cin_out_V_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper257_U0_fifo_cin_out_V_V_din_pass_1_q0 <= PE_wrapper257_U0_fifo_cin_out_V_V_din_pass_1_out;
  end
  assign PE_wrapper257_U0_fifo_cin_out_V_V_din_pass_1_in = PE_wrapper257_U0_fifo_cin_out_V_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_9_11_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_9_11_V_V_full_n_pass_0_q0 <= fifo_cin_PE_9_11_V_V_full_n_pass_0_out;
  end
  assign fifo_cin_PE_9_11_V_V_full_n_pass_0_in = fifo_cin_PE_9_11_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper257_U0_fifo_cin_out_V_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper257_U0_fifo_cin_out_V_V_write_pass_1_q0 <= PE_wrapper257_U0_fifo_cin_out_V_V_write_pass_1_out;
  end
  assign PE_wrapper257_U0_fifo_cin_out_V_V_write_pass_1_in = PE_wrapper257_U0_fifo_cin_out_V_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [63:0] cout_drain_IO_L1_out_wrapper551_U0_fifo_cout_drain_out_V_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper551_U0_fifo_cout_drain_out_V_V_din_pass_1_q0 <= cout_drain_IO_L1_out_wrapper551_U0_fifo_cout_drain_out_V_V_din_pass_1_out;
  end
  assign cout_drain_IO_L1_out_wrapper551_U0_fifo_cout_drain_out_V_V_din_pass_1_in = cout_drain_IO_L1_out_wrapper551_U0_fifo_cout_drain_out_V_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_cout_drain_IO_L1_out_11_6_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_cout_drain_IO_L1_out_11_6_V_V_full_n_pass_0_q0 <= fifo_cout_drain_cout_drain_IO_L1_out_11_6_V_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_cout_drain_IO_L1_out_11_6_V_V_full_n_pass_0_in = fifo_cout_drain_cout_drain_IO_L1_out_11_6_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  cout_drain_IO_L1_out_wrapper551_U0_fifo_cout_drain_out_V_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper551_U0_fifo_cout_drain_out_V_V_write_pass_1_q0 <= cout_drain_IO_L1_out_wrapper551_U0_fifo_cout_drain_out_V_V_write_pass_1_out;
  end
  assign cout_drain_IO_L1_out_wrapper551_U0_fifo_cout_drain_out_V_V_write_pass_1_in = cout_drain_IO_L1_out_wrapper551_U0_fifo_cout_drain_out_V_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper161_U0_fifo_cin_out_V_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper161_U0_fifo_cin_out_V_V_din_pass_1_q0 <= PE_wrapper161_U0_fifo_cin_out_V_V_din_pass_1_out;
  end
  assign PE_wrapper161_U0_fifo_cin_out_V_V_din_pass_1_in = PE_wrapper161_U0_fifo_cin_out_V_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_1_11_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_1_11_V_V_full_n_pass_0_q0 <= fifo_cin_PE_1_11_V_V_full_n_pass_0_out;
  end
  assign fifo_cin_PE_1_11_V_V_full_n_pass_0_in = fifo_cin_PE_1_11_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper161_U0_fifo_cin_out_V_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper161_U0_fifo_cin_out_V_V_write_pass_1_q0 <= PE_wrapper161_U0_fifo_cin_out_V_V_write_pass_1_out;
  end
  assign PE_wrapper161_U0_fifo_cin_out_V_V_write_pass_1_in = PE_wrapper161_U0_fifo_cin_out_V_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [31:0] PE_wrapper185_U0_fifo_cout_drain_out_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper185_U0_fifo_cout_drain_out_V_din_pass_1_q0 <= PE_wrapper185_U0_fifo_cout_drain_out_V_din_pass_1_out;
  end
  assign PE_wrapper185_U0_fifo_cout_drain_out_V_din_pass_1_in = PE_wrapper185_U0_fifo_cout_drain_out_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_PE_2_11_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_PE_2_11_V_full_n_pass_0_q0 <= fifo_cout_drain_PE_2_11_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_PE_2_11_V_full_n_pass_0_in = fifo_cout_drain_PE_2_11_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper185_U0_fifo_cout_drain_out_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper185_U0_fifo_cout_drain_out_V_write_pass_1_q0 <= PE_wrapper185_U0_fifo_cout_drain_out_V_write_pass_1_out;
  end
  assign PE_wrapper185_U0_fifo_cout_drain_out_V_write_pass_1_in = PE_wrapper185_U0_fifo_cout_drain_out_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [63:0] cout_drain_IO_L1_out_wrapper518_U0_fifo_cout_drain_out_V_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper518_U0_fifo_cout_drain_out_V_V_din_pass_1_q0 <= cout_drain_IO_L1_out_wrapper518_U0_fifo_cout_drain_out_V_V_din_pass_1_out;
  end
  assign cout_drain_IO_L1_out_wrapper518_U0_fifo_cout_drain_out_V_V_din_pass_1_in = cout_drain_IO_L1_out_wrapper518_U0_fifo_cout_drain_out_V_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_cout_drain_IO_L1_out_9_8_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_cout_drain_IO_L1_out_9_8_V_V_full_n_pass_0_q0 <= fifo_cout_drain_cout_drain_IO_L1_out_9_8_V_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_cout_drain_IO_L1_out_9_8_V_V_full_n_pass_0_in = fifo_cout_drain_cout_drain_IO_L1_out_9_8_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  cout_drain_IO_L1_out_wrapper518_U0_fifo_cout_drain_out_V_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper518_U0_fifo_cout_drain_out_V_V_write_pass_1_q0 <= cout_drain_IO_L1_out_wrapper518_U0_fifo_cout_drain_out_V_V_write_pass_1_out;
  end
  assign cout_drain_IO_L1_out_wrapper518_U0_fifo_cout_drain_out_V_V_write_pass_1_in = cout_drain_IO_L1_out_wrapper518_U0_fifo_cout_drain_out_V_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [63:0] cout_drain_IO_L1_out_wrapper534_U0_fifo_cout_drain_out_V_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper534_U0_fifo_cout_drain_out_V_V_din_pass_1_q0 <= cout_drain_IO_L1_out_wrapper534_U0_fifo_cout_drain_out_V_V_din_pass_1_out;
  end
  assign cout_drain_IO_L1_out_wrapper534_U0_fifo_cout_drain_out_V_V_din_pass_1_in = cout_drain_IO_L1_out_wrapper534_U0_fifo_cout_drain_out_V_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_cout_drain_IO_L1_out_10_8_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_cout_drain_IO_L1_out_10_8_V_V_full_n_pass_0_q0 <= fifo_cout_drain_cout_drain_IO_L1_out_10_8_V_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_cout_drain_IO_L1_out_10_8_V_V_full_n_pass_0_in = fifo_cout_drain_cout_drain_IO_L1_out_10_8_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  cout_drain_IO_L1_out_wrapper534_U0_fifo_cout_drain_out_V_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper534_U0_fifo_cout_drain_out_V_V_write_pass_1_q0 <= cout_drain_IO_L1_out_wrapper534_U0_fifo_cout_drain_out_V_V_write_pass_1_out;
  end
  assign cout_drain_IO_L1_out_wrapper534_U0_fifo_cout_drain_out_V_V_write_pass_1_in = cout_drain_IO_L1_out_wrapper534_U0_fifo_cout_drain_out_V_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [31:0] PE_wrapper197_U0_fifo_cout_drain_out_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper197_U0_fifo_cout_drain_out_V_din_pass_1_q0 <= PE_wrapper197_U0_fifo_cout_drain_out_V_din_pass_1_out;
  end
  assign PE_wrapper197_U0_fifo_cout_drain_out_V_din_pass_1_in = PE_wrapper197_U0_fifo_cout_drain_out_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_PE_3_11_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_PE_3_11_V_full_n_pass_0_q0 <= fifo_cout_drain_PE_3_11_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_PE_3_11_V_full_n_pass_0_in = fifo_cout_drain_PE_3_11_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper197_U0_fifo_cout_drain_out_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper197_U0_fifo_cout_drain_out_V_write_pass_1_q0 <= PE_wrapper197_U0_fifo_cout_drain_out_V_write_pass_1_out;
  end
  assign PE_wrapper197_U0_fifo_cout_drain_out_V_write_pass_1_in = PE_wrapper197_U0_fifo_cout_drain_out_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [63:0] cout_drain_IO_L1_out_wrapper523_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper523_U0_fifo_cout_drain_out_V_V_din_pass_0_q0 <= cout_drain_IO_L1_out_wrapper523_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper523_U0_fifo_cout_drain_out_V_V_din_pass_0_in = cout_drain_IO_L1_out_wrapper523_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  cout_drain_IO_L1_out_wrapper523_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper523_U0_fifo_cout_drain_out_V_V_write_pass_0_q0 <= cout_drain_IO_L1_out_wrapper523_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper523_U0_fifo_cout_drain_out_V_V_write_pass_0_in = cout_drain_IO_L1_out_wrapper523_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_cout_drain_IO_L1_out_10_7_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_cout_drain_IO_L1_out_10_7_V_V_full_n_pass_0_q0 <= fifo_cout_drain_cout_drain_IO_L1_out_10_7_V_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_cout_drain_IO_L1_out_10_7_V_V_full_n_pass_0_in = fifo_cout_drain_cout_drain_IO_L1_out_10_7_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_cout_drain_IO_L1_out_10_5_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_cout_drain_IO_L1_out_10_5_V_V_full_n_pass_0_q0 <= fifo_cout_drain_cout_drain_IO_L1_out_10_5_V_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_cout_drain_IO_L1_out_10_5_V_V_full_n_pass_0_in = fifo_cout_drain_cout_drain_IO_L1_out_10_5_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_cout_drain_IO_L1_out_11_2_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_cout_drain_IO_L1_out_11_2_V_V_full_n_pass_0_q0 <= fifo_cout_drain_cout_drain_IO_L1_out_11_2_V_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_cout_drain_IO_L1_out_11_2_V_V_full_n_pass_0_in = fifo_cout_drain_cout_drain_IO_L1_out_11_2_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper196_U0_fifo_cin_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper196_U0_fifo_cin_out_V_V_din_pass_0_q0 <= PE_wrapper196_U0_fifo_cin_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper196_U0_fifo_cin_out_V_V_din_pass_0_in = PE_wrapper196_U0_fifo_cin_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper196_U0_fifo_cin_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper196_U0_fifo_cin_out_V_V_write_pass_0_q0 <= PE_wrapper196_U0_fifo_cin_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper196_U0_fifo_cin_out_V_V_write_pass_0_in = PE_wrapper196_U0_fifo_cin_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [63:0] cout_drain_IO_L1_out_wrapper556_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper556_U0_fifo_cout_drain_out_V_V_din_pass_0_q0 <= cout_drain_IO_L1_out_wrapper556_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper556_U0_fifo_cout_drain_out_V_V_din_pass_0_in = cout_drain_IO_L1_out_wrapper556_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  cout_drain_IO_L1_out_wrapper556_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper556_U0_fifo_cout_drain_out_V_V_write_pass_0_q0 <= cout_drain_IO_L1_out_wrapper556_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper556_U0_fifo_cout_drain_out_V_V_write_pass_0_in = cout_drain_IO_L1_out_wrapper556_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [63:0] cout_drain_IO_L1_out_wrapper539_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper539_U0_fifo_cout_drain_out_V_V_din_pass_0_q0 <= cout_drain_IO_L1_out_wrapper539_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper539_U0_fifo_cout_drain_out_V_V_din_pass_0_in = cout_drain_IO_L1_out_wrapper539_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  cout_drain_IO_L1_out_wrapper539_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper539_U0_fifo_cout_drain_out_V_V_write_pass_0_q0 <= cout_drain_IO_L1_out_wrapper539_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper539_U0_fifo_cout_drain_out_V_V_write_pass_0_in = cout_drain_IO_L1_out_wrapper539_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper231_U0_fifo_w_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper231_U0_fifo_w_out_V_V_din_pass_0_q0 <= PE_wrapper231_U0_fifo_w_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper231_U0_fifo_w_out_V_V_din_pass_0_in = PE_wrapper231_U0_fifo_w_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper231_U0_fifo_w_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper231_U0_fifo_w_out_V_V_write_pass_0_q0 <= PE_wrapper231_U0_fifo_w_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper231_U0_fifo_w_out_V_V_write_pass_0_in = PE_wrapper231_U0_fifo_w_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [31:0] PE_wrapper231_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper231_U0_fifo_cout_drain_out_V_din_pass_0_q0 <= PE_wrapper231_U0_fifo_cout_drain_out_V_din_pass_0_out;
  end
  assign PE_wrapper231_U0_fifo_cout_drain_out_V_din_pass_0_in = PE_wrapper231_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper231_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper231_U0_fifo_cout_drain_out_V_write_pass_0_q0 <= PE_wrapper231_U0_fifo_cout_drain_out_V_write_pass_0_out;
  end
  assign PE_wrapper231_U0_fifo_cout_drain_out_V_write_pass_0_in = PE_wrapper231_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_6_9_V_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_6_9_V_V_full_n_pass_1_q0 <= fifo_w_PE_6_9_V_V_full_n_pass_1_out;
  end
  assign fifo_w_PE_6_9_V_V_full_n_pass_1_in = fifo_w_PE_6_9_V_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg [63:0] cout_drain_IO_L2_out558_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L2_out558_U0_fifo_cout_drain_out_V_V_din_pass_0_q0 <= cout_drain_IO_L2_out558_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  end
  assign cout_drain_IO_L2_out558_U0_fifo_cout_drain_out_V_V_din_pass_0_in = cout_drain_IO_L2_out558_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  cout_drain_IO_L2_out558_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L2_out558_U0_fifo_cout_drain_out_V_V_write_pass_0_q0 <= cout_drain_IO_L2_out558_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  end
  assign cout_drain_IO_L2_out558_U0_fifo_cout_drain_out_V_V_write_pass_0_in = cout_drain_IO_L2_out558_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [31:0] PE_wrapper221_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper221_U0_fifo_cout_drain_out_V_din_pass_0_q0 <= PE_wrapper221_U0_fifo_cout_drain_out_V_din_pass_0_out;
  end
  assign PE_wrapper221_U0_fifo_cout_drain_out_V_din_pass_0_in = PE_wrapper221_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper221_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper221_U0_fifo_cout_drain_out_V_write_pass_0_q0 <= PE_wrapper221_U0_fifo_cout_drain_out_V_write_pass_0_out;
  end
  assign PE_wrapper221_U0_fifo_cout_drain_out_V_write_pass_0_in = PE_wrapper221_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper184_U0_fifo_w_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper184_U0_fifo_w_out_V_V_din_pass_0_q0 <= PE_wrapper184_U0_fifo_w_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper184_U0_fifo_w_out_V_V_din_pass_0_in = PE_wrapper184_U0_fifo_w_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper184_U0_fifo_w_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper184_U0_fifo_w_out_V_V_write_pass_0_q0 <= PE_wrapper184_U0_fifo_w_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper184_U0_fifo_w_out_V_V_write_pass_0_in = PE_wrapper184_U0_fifo_w_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_PE_6_10_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_PE_6_10_V_full_n_pass_0_q0 <= fifo_cout_drain_PE_6_10_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_PE_6_10_V_full_n_pass_0_in = fifo_cout_drain_PE_6_10_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_cout_drain_IO_L1_out_9_4_V_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_cout_drain_IO_L1_out_9_4_V_V_full_n_pass_1_q0 <= fifo_cout_drain_cout_drain_IO_L1_out_9_4_V_V_full_n_pass_1_out;
  end
  assign fifo_cout_drain_cout_drain_IO_L1_out_9_4_V_V_full_n_pass_1_in = fifo_cout_drain_cout_drain_IO_L1_out_9_4_V_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper196_U0_fifo_w_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper196_U0_fifo_w_out_V_V_din_pass_0_q0 <= PE_wrapper196_U0_fifo_w_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper196_U0_fifo_w_out_V_V_din_pass_0_in = PE_wrapper196_U0_fifo_w_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper196_U0_fifo_w_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper196_U0_fifo_w_out_V_V_write_pass_0_q0 <= PE_wrapper196_U0_fifo_w_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper196_U0_fifo_w_out_V_V_write_pass_0_in = PE_wrapper196_U0_fifo_w_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper209_U0_fifo_w_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper209_U0_fifo_w_out_V_V_din_pass_0_q0 <= PE_wrapper209_U0_fifo_w_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper209_U0_fifo_w_out_V_V_din_pass_0_in = PE_wrapper209_U0_fifo_w_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper209_U0_fifo_w_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper209_U0_fifo_w_out_V_V_write_pass_0_q0 <= PE_wrapper209_U0_fifo_w_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper209_U0_fifo_w_out_V_V_write_pass_0_in = PE_wrapper209_U0_fifo_w_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_cout_drain_IO_L1_out_11_5_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_cout_drain_IO_L1_out_11_5_V_V_full_n_pass_0_q0 <= fifo_cout_drain_cout_drain_IO_L1_out_11_5_V_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_cout_drain_IO_L1_out_11_5_V_V_full_n_pass_0_in = fifo_cout_drain_cout_drain_IO_L1_out_11_5_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper233_U0_fifo_cin_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper233_U0_fifo_cin_out_V_V_din_pass_0_q0 <= PE_wrapper233_U0_fifo_cin_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper233_U0_fifo_cin_out_V_V_din_pass_0_in = PE_wrapper233_U0_fifo_cin_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper233_U0_fifo_cin_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper233_U0_fifo_cin_out_V_V_write_pass_0_q0 <= PE_wrapper233_U0_fifo_cin_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper233_U0_fifo_cin_out_V_V_write_pass_0_in = PE_wrapper233_U0_fifo_cin_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [31:0] PE_wrapper184_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper184_U0_fifo_cout_drain_out_V_din_pass_0_q0 <= PE_wrapper184_U0_fifo_cout_drain_out_V_din_pass_0_out;
  end
  assign PE_wrapper184_U0_fifo_cout_drain_out_V_din_pass_0_in = PE_wrapper184_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper184_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper184_U0_fifo_cout_drain_out_V_write_pass_0_q0 <= PE_wrapper184_U0_fifo_cout_drain_out_V_write_pass_0_out;
  end
  assign PE_wrapper184_U0_fifo_cout_drain_out_V_write_pass_0_in = PE_wrapper184_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_cout_drain_IO_L2_out_11_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_cout_drain_IO_L2_out_11_V_V_full_n_pass_0_q0 <= fifo_cout_drain_cout_drain_IO_L2_out_11_V_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_cout_drain_IO_L2_out_11_V_V_full_n_pass_0_in = fifo_cout_drain_cout_drain_IO_L2_out_11_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_4_11_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_4_11_V_V_full_n_pass_0_q0 <= fifo_cin_PE_4_11_V_V_full_n_pass_0_out;
  end
  assign fifo_cin_PE_4_11_V_V_full_n_pass_0_in = fifo_cin_PE_4_11_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_cout_drain_IO_L1_out_10_0_V_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_cout_drain_IO_L1_out_10_0_V_V_full_n_pass_1_q0 <= fifo_cout_drain_cout_drain_IO_L1_out_10_0_V_V_full_n_pass_1_out;
  end
  assign fifo_cout_drain_cout_drain_IO_L1_out_10_0_V_V_full_n_pass_1_in = fifo_cout_drain_cout_drain_IO_L1_out_10_0_V_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_6_9_V_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_6_9_V_V_full_n_pass_1_q0 <= fifo_cin_PE_6_9_V_V_full_n_pass_1_out;
  end
  assign fifo_cin_PE_6_9_V_V_full_n_pass_1_in = fifo_cin_PE_6_9_V_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_PE_1_11_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_PE_1_11_V_full_n_pass_0_q0 <= fifo_cout_drain_PE_1_11_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_PE_1_11_V_full_n_pass_0_in = fifo_cout_drain_PE_1_11_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg [63:0] cout_drain_IO_L1_out_wrapper549_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper549_U0_fifo_cout_drain_out_V_V_din_pass_0_q0 <= cout_drain_IO_L1_out_wrapper549_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper549_U0_fifo_cout_drain_out_V_V_din_pass_0_in = cout_drain_IO_L1_out_wrapper549_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  cout_drain_IO_L1_out_wrapper549_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper549_U0_fifo_cout_drain_out_V_V_write_pass_0_q0 <= cout_drain_IO_L1_out_wrapper549_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper549_U0_fifo_cout_drain_out_V_V_write_pass_0_in = cout_drain_IO_L1_out_wrapper549_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_2_10_V_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_2_10_V_V_full_n_pass_1_q0 <= fifo_cin_PE_2_10_V_V_full_n_pass_1_out;
  end
  assign fifo_cin_PE_2_10_V_V_full_n_pass_1_in = fifo_cin_PE_2_10_V_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper195_U0_fifo_cin_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper195_U0_fifo_cin_out_V_V_din_pass_0_q0 <= PE_wrapper195_U0_fifo_cin_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper195_U0_fifo_cin_out_V_V_din_pass_0_in = PE_wrapper195_U0_fifo_cin_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper195_U0_fifo_cin_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper195_U0_fifo_cin_out_V_V_write_pass_0_q0 <= PE_wrapper195_U0_fifo_cin_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper195_U0_fifo_cin_out_V_V_write_pass_0_in = PE_wrapper195_U0_fifo_cin_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [63:0] cout_drain_IO_L1_out_wrapper536_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper536_U0_fifo_cout_drain_out_V_V_din_pass_0_q0 <= cout_drain_IO_L1_out_wrapper536_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper536_U0_fifo_cout_drain_out_V_V_din_pass_0_in = cout_drain_IO_L1_out_wrapper536_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  cout_drain_IO_L1_out_wrapper536_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper536_U0_fifo_cout_drain_out_V_V_write_pass_0_q0 <= cout_drain_IO_L1_out_wrapper536_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper536_U0_fifo_cout_drain_out_V_V_write_pass_0_in = cout_drain_IO_L1_out_wrapper536_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_PE_4_10_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_PE_4_10_V_full_n_pass_0_q0 <= fifo_cout_drain_PE_4_10_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_PE_4_10_V_full_n_pass_0_in = fifo_cout_drain_PE_4_10_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_5_11_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_5_11_V_V_full_n_pass_0_q0 <= fifo_w_PE_5_11_V_V_full_n_pass_0_out;
  end
  assign fifo_w_PE_5_11_V_V_full_n_pass_0_in = fifo_w_PE_5_11_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_cin_IO_L2_in_11_V_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_cin_IO_L2_in_11_V_V_full_n_pass_1_q0 <= fifo_cin_cin_IO_L2_in_11_V_V_full_n_pass_1_out;
  end
  assign fifo_cin_cin_IO_L2_in_11_V_V_full_n_pass_1_in = fifo_cin_cin_IO_L2_in_11_V_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_cout_drain_IO_L1_out_9_6_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_cout_drain_IO_L1_out_9_6_V_V_full_n_pass_0_q0 <= fifo_cout_drain_cout_drain_IO_L1_out_9_6_V_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_cout_drain_IO_L1_out_9_6_V_V_full_n_pass_0_in = fifo_cout_drain_cout_drain_IO_L1_out_9_6_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_PE_8_11_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_PE_8_11_V_full_n_pass_0_q0 <= fifo_cout_drain_PE_8_11_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_PE_8_11_V_full_n_pass_0_in = fifo_cout_drain_PE_8_11_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] cin_IO_L2_in_boundary_U0_fifo_cin_local_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    cin_IO_L2_in_boundary_U0_fifo_cin_local_out_V_V_din_pass_0_q0 <= cin_IO_L2_in_boundary_U0_fifo_cin_local_out_V_V_din_pass_0_out;
  end
  assign cin_IO_L2_in_boundary_U0_fifo_cin_local_out_V_V_din_pass_0_in = cin_IO_L2_in_boundary_U0_fifo_cin_local_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  cin_IO_L2_in_boundary_U0_fifo_cin_local_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    cin_IO_L2_in_boundary_U0_fifo_cin_local_out_V_V_write_pass_0_q0 <= cin_IO_L2_in_boundary_U0_fifo_cin_local_out_V_V_write_pass_0_out;
  end
  assign cin_IO_L2_in_boundary_U0_fifo_cin_local_out_V_V_write_pass_0_in = cin_IO_L2_in_boundary_U0_fifo_cin_local_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_6_11_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_6_11_V_V_full_n_pass_0_q0 <= fifo_w_PE_6_11_V_V_full_n_pass_0_out;
  end
  assign fifo_w_PE_6_11_V_V_full_n_pass_0_in = fifo_w_PE_6_11_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_2_10_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_2_10_V_V_full_n_pass_0_q0 <= fifo_w_PE_2_10_V_V_full_n_pass_0_out;
  end
  assign fifo_w_PE_2_10_V_V_full_n_pass_0_in = fifo_w_PE_2_10_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper221_U0_fifo_w_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper221_U0_fifo_w_out_V_V_din_pass_0_q0 <= PE_wrapper221_U0_fifo_w_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper221_U0_fifo_w_out_V_V_din_pass_0_in = PE_wrapper221_U0_fifo_w_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper221_U0_fifo_w_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper221_U0_fifo_w_out_V_V_write_pass_0_q0 <= PE_wrapper221_U0_fifo_w_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper221_U0_fifo_w_out_V_V_write_pass_0_in = PE_wrapper221_U0_fifo_w_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_4_11_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_4_11_V_V_full_n_pass_0_q0 <= fifo_w_PE_4_11_V_V_full_n_pass_0_out;
  end
  assign fifo_w_PE_4_11_V_V_full_n_pass_0_in = fifo_w_PE_4_11_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg [31:0] PE_wrapper233_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper233_U0_fifo_cout_drain_out_V_din_pass_0_q0 <= PE_wrapper233_U0_fifo_cout_drain_out_V_din_pass_0_out;
  end
  assign PE_wrapper233_U0_fifo_cout_drain_out_V_din_pass_0_in = PE_wrapper233_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper233_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper233_U0_fifo_cout_drain_out_V_write_pass_0_q0 <= PE_wrapper233_U0_fifo_cout_drain_out_V_write_pass_0_out;
  end
  assign PE_wrapper233_U0_fifo_cout_drain_out_V_write_pass_0_in = PE_wrapper233_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_3_9_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_3_9_V_V_full_n_pass_0_q0 <= fifo_cin_PE_3_9_V_V_full_n_pass_0_out;
  end
  assign fifo_cin_PE_3_9_V_V_full_n_pass_0_in = fifo_cin_PE_3_9_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_3_9_V_V_full_n_pass_2_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_3_9_V_V_full_n_pass_2_q0 <= fifo_w_PE_3_9_V_V_full_n_pass_2_out;
  end
  assign fifo_w_PE_3_9_V_V_full_n_pass_2_in = fifo_w_PE_3_9_V_V_full_n_pass_2_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper231_U0_fifo_cin_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper231_U0_fifo_cin_out_V_V_din_pass_0_q0 <= PE_wrapper231_U0_fifo_cin_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper231_U0_fifo_cin_out_V_V_din_pass_0_in = PE_wrapper231_U0_fifo_cin_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper231_U0_fifo_cin_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper231_U0_fifo_cin_out_V_V_write_pass_0_q0 <= PE_wrapper231_U0_fifo_cin_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper231_U0_fifo_cin_out_V_V_write_pass_0_in = PE_wrapper231_U0_fifo_cin_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_2_12_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_2_12_V_V_full_n_pass_0_q0 <= fifo_w_PE_2_12_V_V_full_n_pass_0_out;
  end
  assign fifo_w_PE_2_12_V_V_full_n_pass_0_in = fifo_w_PE_2_12_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_cout_drain_IO_L1_out_11_9_V_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_cout_drain_IO_L1_out_11_9_V_V_full_n_pass_1_q0 <= fifo_cout_drain_cout_drain_IO_L1_out_11_9_V_V_full_n_pass_1_out;
  end
  assign fifo_cout_drain_cout_drain_IO_L1_out_11_9_V_V_full_n_pass_1_in = fifo_cout_drain_cout_drain_IO_L1_out_11_9_V_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg [63:0] cout_drain_IO_L1_out_wrapper521_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper521_U0_fifo_cout_drain_out_V_V_din_pass_0_q0 <= cout_drain_IO_L1_out_wrapper521_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper521_U0_fifo_cout_drain_out_V_V_din_pass_0_in = cout_drain_IO_L1_out_wrapper521_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  cout_drain_IO_L1_out_wrapper521_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper521_U0_fifo_cout_drain_out_V_V_write_pass_0_q0 <= cout_drain_IO_L1_out_wrapper521_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper521_U0_fifo_cout_drain_out_V_V_write_pass_0_in = cout_drain_IO_L1_out_wrapper521_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_PE_5_9_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_PE_5_9_V_full_n_pass_1_q0 <= fifo_cout_drain_PE_5_9_V_full_n_pass_1_out;
  end
  assign fifo_cout_drain_PE_5_9_V_full_n_pass_1_in = fifo_cout_drain_PE_5_9_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg [63:0] cout_drain_IO_L1_out_wrapper553_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper553_U0_fifo_cout_drain_out_V_V_din_pass_0_q0 <= cout_drain_IO_L1_out_wrapper553_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper553_U0_fifo_cout_drain_out_V_V_din_pass_0_in = cout_drain_IO_L1_out_wrapper553_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  cout_drain_IO_L1_out_wrapper553_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper553_U0_fifo_cout_drain_out_V_V_write_pass_0_q0 <= cout_drain_IO_L1_out_wrapper553_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper553_U0_fifo_cout_drain_out_V_V_write_pass_0_in = cout_drain_IO_L1_out_wrapper553_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  ap_done_Boundary_X4Y14_To_X6Y14_q0;
  always @ (posedge ap_clk) begin
    ap_done_Boundary_X4Y14_To_X6Y14_q0 <= ap_done_Boundary_X4Y14_To_X6Y14_out;
  end
  assign ap_done_Boundary_X4Y14_To_X6Y14_in = ap_done_Boundary_X4Y14_To_X6Y14_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper231_U0_fifo_cin_out_V_V_din_pass_2_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper231_U0_fifo_cin_out_V_V_din_pass_2_q0 <= PE_wrapper231_U0_fifo_cin_out_V_V_din_pass_2_out;
  end
  assign PE_wrapper231_U0_fifo_cin_out_V_V_din_pass_2_in = PE_wrapper231_U0_fifo_cin_out_V_V_din_pass_2_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_7_9_V_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_7_9_V_V_full_n_pass_1_q0 <= fifo_cin_PE_7_9_V_V_full_n_pass_1_out;
  end
  assign fifo_cin_PE_7_9_V_V_full_n_pass_1_in = fifo_cin_PE_7_9_V_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper231_U0_fifo_cin_out_V_V_write_pass_2_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper231_U0_fifo_cin_out_V_V_write_pass_2_q0 <= PE_wrapper231_U0_fifo_cin_out_V_V_write_pass_2_out;
  end
  assign PE_wrapper231_U0_fifo_cin_out_V_V_write_pass_2_in = PE_wrapper231_U0_fifo_cin_out_V_V_write_pass_2_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper244_U0_fifo_cin_out_V_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper244_U0_fifo_cin_out_V_V_din_pass_1_q0 <= PE_wrapper244_U0_fifo_cin_out_V_V_din_pass_1_out;
  end
  assign PE_wrapper244_U0_fifo_cin_out_V_V_din_pass_1_in = PE_wrapper244_U0_fifo_cin_out_V_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_8_10_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_8_10_V_V_full_n_pass_0_q0 <= fifo_cin_PE_8_10_V_V_full_n_pass_0_out;
  end
  assign fifo_cin_PE_8_10_V_V_full_n_pass_0_in = fifo_cin_PE_8_10_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper244_U0_fifo_cin_out_V_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper244_U0_fifo_cin_out_V_V_write_pass_1_q0 <= PE_wrapper244_U0_fifo_cin_out_V_V_write_pass_1_out;
  end
  assign PE_wrapper244_U0_fifo_cin_out_V_V_write_pass_1_in = PE_wrapper244_U0_fifo_cin_out_V_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper173_U0_fifo_w_out_V_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper173_U0_fifo_w_out_V_V_din_pass_1_q0 <= PE_wrapper173_U0_fifo_w_out_V_V_din_pass_1_out;
  end
  assign PE_wrapper173_U0_fifo_w_out_V_V_din_pass_1_in = PE_wrapper173_U0_fifo_w_out_V_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_1_12_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_1_12_V_V_full_n_pass_0_q0 <= fifo_w_PE_1_12_V_V_full_n_pass_0_out;
  end
  assign fifo_w_PE_1_12_V_V_full_n_pass_0_in = fifo_w_PE_1_12_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper173_U0_fifo_w_out_V_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper173_U0_fifo_w_out_V_V_write_pass_1_q0 <= PE_wrapper173_U0_fifo_w_out_V_V_write_pass_1_out;
  end
  assign PE_wrapper173_U0_fifo_w_out_V_V_write_pass_1_in = PE_wrapper173_U0_fifo_w_out_V_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [31:0] PE_wrapper255_U0_fifo_cout_drain_out_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper255_U0_fifo_cout_drain_out_V_din_pass_1_q0 <= PE_wrapper255_U0_fifo_cout_drain_out_V_din_pass_1_out;
  end
  assign PE_wrapper255_U0_fifo_cout_drain_out_V_din_pass_1_in = PE_wrapper255_U0_fifo_cout_drain_out_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_PE_8_9_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_PE_8_9_V_full_n_pass_0_q0 <= fifo_cout_drain_PE_8_9_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_PE_8_9_V_full_n_pass_0_in = fifo_cout_drain_PE_8_9_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper255_U0_fifo_cout_drain_out_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper255_U0_fifo_cout_drain_out_V_write_pass_1_q0 <= PE_wrapper255_U0_fifo_cout_drain_out_V_write_pass_1_out;
  end
  assign PE_wrapper255_U0_fifo_cout_drain_out_V_write_pass_1_in = PE_wrapper255_U0_fifo_cout_drain_out_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper244_U0_fifo_w_out_V_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper244_U0_fifo_w_out_V_V_din_pass_1_q0 <= PE_wrapper244_U0_fifo_w_out_V_V_din_pass_1_out;
  end
  assign PE_wrapper244_U0_fifo_w_out_V_V_din_pass_1_in = PE_wrapper244_U0_fifo_w_out_V_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_7_11_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_7_11_V_V_full_n_pass_0_q0 <= fifo_w_PE_7_11_V_V_full_n_pass_0_out;
  end
  assign fifo_w_PE_7_11_V_V_full_n_pass_0_in = fifo_w_PE_7_11_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper244_U0_fifo_w_out_V_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper244_U0_fifo_w_out_V_V_write_pass_1_q0 <= PE_wrapper244_U0_fifo_w_out_V_V_write_pass_1_out;
  end
  assign PE_wrapper244_U0_fifo_w_out_V_V_write_pass_1_in = PE_wrapper244_U0_fifo_w_out_V_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [63:0] cout_drain_IO_L1_out_wrapper517_U0_fifo_cout_drain_out_V_V_din_pass_2_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper517_U0_fifo_cout_drain_out_V_V_din_pass_2_q0 <= cout_drain_IO_L1_out_wrapper517_U0_fifo_cout_drain_out_V_V_din_pass_2_out;
  end
  assign cout_drain_IO_L1_out_wrapper517_U0_fifo_cout_drain_out_V_V_din_pass_2_in = cout_drain_IO_L1_out_wrapper517_U0_fifo_cout_drain_out_V_V_din_pass_2_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_cout_drain_IO_L1_out_9_9_V_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_cout_drain_IO_L1_out_9_9_V_V_full_n_pass_1_q0 <= fifo_cout_drain_cout_drain_IO_L1_out_9_9_V_V_full_n_pass_1_out;
  end
  assign fifo_cout_drain_cout_drain_IO_L1_out_9_9_V_V_full_n_pass_1_in = fifo_cout_drain_cout_drain_IO_L1_out_9_9_V_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg  cout_drain_IO_L1_out_wrapper517_U0_fifo_cout_drain_out_V_V_write_pass_2_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper517_U0_fifo_cout_drain_out_V_V_write_pass_2_q0 <= cout_drain_IO_L1_out_wrapper517_U0_fifo_cout_drain_out_V_V_write_pass_2_out;
  end
  assign cout_drain_IO_L1_out_wrapper517_U0_fifo_cout_drain_out_V_V_write_pass_2_in = cout_drain_IO_L1_out_wrapper517_U0_fifo_cout_drain_out_V_V_write_pass_2_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper255_U0_fifo_w_out_V_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper255_U0_fifo_w_out_V_V_din_pass_1_q0 <= PE_wrapper255_U0_fifo_w_out_V_V_din_pass_1_out;
  end
  assign PE_wrapper255_U0_fifo_w_out_V_V_din_pass_1_in = PE_wrapper255_U0_fifo_w_out_V_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_8_10_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_8_10_V_V_full_n_pass_0_q0 <= fifo_w_PE_8_10_V_V_full_n_pass_0_out;
  end
  assign fifo_w_PE_8_10_V_V_full_n_pass_0_in = fifo_w_PE_8_10_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper255_U0_fifo_w_out_V_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper255_U0_fifo_w_out_V_V_write_pass_1_q0 <= PE_wrapper255_U0_fifo_w_out_V_V_write_pass_1_out;
  end
  assign PE_wrapper255_U0_fifo_w_out_V_V_write_pass_1_in = PE_wrapper255_U0_fifo_w_out_V_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper173_U0_fifo_cin_out_V_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper173_U0_fifo_cin_out_V_V_din_pass_1_q0 <= PE_wrapper173_U0_fifo_cin_out_V_V_din_pass_1_out;
  end
  assign PE_wrapper173_U0_fifo_cin_out_V_V_din_pass_1_in = PE_wrapper173_U0_fifo_cin_out_V_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_2_11_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_2_11_V_V_full_n_pass_0_q0 <= fifo_cin_PE_2_11_V_V_full_n_pass_0_out;
  end
  assign fifo_cin_PE_2_11_V_V_full_n_pass_0_in = fifo_cin_PE_2_11_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper173_U0_fifo_cin_out_V_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper173_U0_fifo_cin_out_V_V_write_pass_1_q0 <= PE_wrapper173_U0_fifo_cin_out_V_V_write_pass_1_out;
  end
  assign PE_wrapper173_U0_fifo_cin_out_V_V_write_pass_1_in = PE_wrapper173_U0_fifo_cin_out_V_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [63:0] cout_drain_IO_L1_out_wrapper533_U0_fifo_cout_drain_out_V_V_din_pass_2_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper533_U0_fifo_cout_drain_out_V_V_din_pass_2_q0 <= cout_drain_IO_L1_out_wrapper533_U0_fifo_cout_drain_out_V_V_din_pass_2_out;
  end
  assign cout_drain_IO_L1_out_wrapper533_U0_fifo_cout_drain_out_V_V_din_pass_2_in = cout_drain_IO_L1_out_wrapper533_U0_fifo_cout_drain_out_V_V_din_pass_2_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_cout_drain_IO_L1_out_10_9_V_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_cout_drain_IO_L1_out_10_9_V_V_full_n_pass_1_q0 <= fifo_cout_drain_cout_drain_IO_L1_out_10_9_V_V_full_n_pass_1_out;
  end
  assign fifo_cout_drain_cout_drain_IO_L1_out_10_9_V_V_full_n_pass_1_in = fifo_cout_drain_cout_drain_IO_L1_out_10_9_V_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg  cout_drain_IO_L1_out_wrapper533_U0_fifo_cout_drain_out_V_V_write_pass_2_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper533_U0_fifo_cout_drain_out_V_V_write_pass_2_q0 <= cout_drain_IO_L1_out_wrapper533_U0_fifo_cout_drain_out_V_V_write_pass_2_out;
  end
  assign cout_drain_IO_L1_out_wrapper533_U0_fifo_cout_drain_out_V_V_write_pass_2_in = cout_drain_IO_L1_out_wrapper533_U0_fifo_cout_drain_out_V_V_write_pass_2_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_0_9_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_0_9_V_V_full_n_pass_0_q0 <= fifo_w_PE_0_9_V_V_full_n_pass_0_out;
  end
  assign fifo_w_PE_0_9_V_V_full_n_pass_0_in = fifo_w_PE_0_9_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_cout_drain_IO_L1_out_9_3_V_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_cout_drain_IO_L1_out_9_3_V_V_full_n_pass_1_q0 <= fifo_cout_drain_cout_drain_IO_L1_out_9_3_V_V_full_n_pass_1_out;
  end
  assign fifo_cout_drain_cout_drain_IO_L1_out_9_3_V_V_full_n_pass_1_in = fifo_cout_drain_cout_drain_IO_L1_out_9_3_V_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper219_U0_fifo_w_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper219_U0_fifo_w_out_V_V_din_pass_0_q0 <= PE_wrapper219_U0_fifo_w_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper219_U0_fifo_w_out_V_V_din_pass_0_in = PE_wrapper219_U0_fifo_w_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper219_U0_fifo_w_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper219_U0_fifo_w_out_V_V_write_pass_0_q0 <= PE_wrapper219_U0_fifo_w_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper219_U0_fifo_w_out_V_V_write_pass_0_in = PE_wrapper219_U0_fifo_w_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_1_9_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_1_9_V_V_full_n_pass_0_q0 <= fifo_w_PE_1_9_V_V_full_n_pass_0_out;
  end
  assign fifo_w_PE_1_9_V_V_full_n_pass_0_in = fifo_w_PE_1_9_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper171_U0_fifo_cin_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper171_U0_fifo_cin_out_V_V_din_pass_0_q0 <= PE_wrapper171_U0_fifo_cin_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper171_U0_fifo_cin_out_V_V_din_pass_0_in = PE_wrapper171_U0_fifo_cin_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper171_U0_fifo_cin_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper171_U0_fifo_cin_out_V_V_write_pass_0_q0 <= PE_wrapper171_U0_fifo_cin_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper171_U0_fifo_cin_out_V_V_write_pass_0_in = PE_wrapper171_U0_fifo_cin_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper172_U0_fifo_w_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper172_U0_fifo_w_out_V_V_din_pass_0_q0 <= PE_wrapper172_U0_fifo_w_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper172_U0_fifo_w_out_V_V_din_pass_0_in = PE_wrapper172_U0_fifo_w_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper172_U0_fifo_w_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper172_U0_fifo_w_out_V_V_write_pass_0_q0 <= PE_wrapper172_U0_fifo_w_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper172_U0_fifo_w_out_V_V_write_pass_0_in = PE_wrapper172_U0_fifo_w_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [63:0] cout_drain_IO_L2_out559_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L2_out559_U0_fifo_cout_drain_out_V_V_din_pass_0_q0 <= cout_drain_IO_L2_out559_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  end
  assign cout_drain_IO_L2_out559_U0_fifo_cout_drain_out_V_V_din_pass_0_in = cout_drain_IO_L2_out559_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  cout_drain_IO_L2_out559_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L2_out559_U0_fifo_cout_drain_out_V_V_write_pass_0_q0 <= cout_drain_IO_L2_out559_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  end
  assign cout_drain_IO_L2_out559_U0_fifo_cout_drain_out_V_V_write_pass_0_in = cout_drain_IO_L2_out559_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_4_9_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_4_9_V_V_full_n_pass_0_q0 <= fifo_w_PE_4_9_V_V_full_n_pass_0_out;
  end
  assign fifo_w_PE_4_9_V_V_full_n_pass_0_in = fifo_w_PE_4_9_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_cin_IO_L2_in_9_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_cin_IO_L2_in_9_V_V_full_n_pass_0_q0 <= fifo_cin_cin_IO_L2_in_9_V_V_full_n_pass_0_out;
  end
  assign fifo_cin_cin_IO_L2_in_9_V_V_full_n_pass_0_in = fifo_cin_cin_IO_L2_in_9_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper160_U0_fifo_w_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper160_U0_fifo_w_out_V_V_din_pass_0_q0 <= PE_wrapper160_U0_fifo_w_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper160_U0_fifo_w_out_V_V_din_pass_0_in = PE_wrapper160_U0_fifo_w_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper160_U0_fifo_w_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper160_U0_fifo_w_out_V_V_write_pass_0_q0 <= PE_wrapper160_U0_fifo_w_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper160_U0_fifo_w_out_V_V_write_pass_0_in = PE_wrapper160_U0_fifo_w_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_cout_drain_IO_L2_out_10_V_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_cout_drain_IO_L2_out_10_V_V_full_n_pass_1_q0 <= fifo_cout_drain_cout_drain_IO_L2_out_10_V_V_full_n_pass_1_out;
  end
  assign fifo_cout_drain_cout_drain_IO_L2_out_10_V_V_full_n_pass_1_in = fifo_cout_drain_cout_drain_IO_L2_out_10_V_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper207_U0_fifo_w_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper207_U0_fifo_w_out_V_V_din_pass_0_q0 <= PE_wrapper207_U0_fifo_w_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper207_U0_fifo_w_out_V_V_din_pass_0_in = PE_wrapper207_U0_fifo_w_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper207_U0_fifo_w_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper207_U0_fifo_w_out_V_V_write_pass_0_q0 <= PE_wrapper207_U0_fifo_w_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper207_U0_fifo_w_out_V_V_write_pass_0_in = PE_wrapper207_U0_fifo_w_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_PE_2_9_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_PE_2_9_V_full_n_pass_0_q0 <= fifo_cout_drain_PE_2_9_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_PE_2_9_V_full_n_pass_0_in = fifo_cout_drain_PE_2_9_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg [63:0] cout_drain_IO_L1_out_wrapper522_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper522_U0_fifo_cout_drain_out_V_V_din_pass_0_q0 <= cout_drain_IO_L1_out_wrapper522_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper522_U0_fifo_cout_drain_out_V_V_din_pass_0_in = cout_drain_IO_L1_out_wrapper522_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  cout_drain_IO_L1_out_wrapper522_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper522_U0_fifo_cout_drain_out_V_V_write_pass_0_q0 <= cout_drain_IO_L1_out_wrapper522_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper522_U0_fifo_cout_drain_out_V_V_write_pass_0_in = cout_drain_IO_L1_out_wrapper522_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_cout_drain_IO_L1_out_10_2_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_cout_drain_IO_L1_out_10_2_V_V_full_n_pass_0_q0 <= fifo_cout_drain_cout_drain_IO_L1_out_10_2_V_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_cout_drain_IO_L1_out_10_2_V_V_full_n_pass_0_in = fifo_cout_drain_cout_drain_IO_L1_out_10_2_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg [63:0] cout_drain_IO_L1_out_wrapper542_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper542_U0_fifo_cout_drain_out_V_V_din_pass_0_q0 <= cout_drain_IO_L1_out_wrapper542_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper542_U0_fifo_cout_drain_out_V_V_din_pass_0_in = cout_drain_IO_L1_out_wrapper542_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  cout_drain_IO_L1_out_wrapper542_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper542_U0_fifo_cout_drain_out_V_V_write_pass_0_q0 <= cout_drain_IO_L1_out_wrapper542_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper542_U0_fifo_cout_drain_out_V_V_write_pass_0_in = cout_drain_IO_L1_out_wrapper542_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper219_U0_fifo_cin_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper219_U0_fifo_cin_out_V_V_din_pass_0_q0 <= PE_wrapper219_U0_fifo_cin_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper219_U0_fifo_cin_out_V_V_din_pass_0_in = PE_wrapper219_U0_fifo_cin_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper219_U0_fifo_cin_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper219_U0_fifo_cin_out_V_V_write_pass_0_q0 <= PE_wrapper219_U0_fifo_cin_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper219_U0_fifo_cin_out_V_V_write_pass_0_in = PE_wrapper219_U0_fifo_cin_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper172_U0_fifo_cin_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper172_U0_fifo_cin_out_V_V_din_pass_0_q0 <= PE_wrapper172_U0_fifo_cin_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper172_U0_fifo_cin_out_V_V_din_pass_0_in = PE_wrapper172_U0_fifo_cin_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper172_U0_fifo_cin_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper172_U0_fifo_cin_out_V_V_write_pass_0_q0 <= PE_wrapper172_U0_fifo_cin_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper172_U0_fifo_cin_out_V_V_write_pass_0_in = PE_wrapper172_U0_fifo_cin_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_4_9_V_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_4_9_V_V_full_n_pass_1_q0 <= fifo_cin_PE_4_9_V_V_full_n_pass_1_out;
  end
  assign fifo_cin_PE_4_9_V_V_full_n_pass_1_in = fifo_cin_PE_4_9_V_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg [255:0] cin_IO_L2_in134_U0_fifo_cin_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    cin_IO_L2_in134_U0_fifo_cin_out_V_V_din_pass_0_q0 <= cin_IO_L2_in134_U0_fifo_cin_out_V_V_din_pass_0_out;
  end
  assign cin_IO_L2_in134_U0_fifo_cin_out_V_V_din_pass_0_in = cin_IO_L2_in134_U0_fifo_cin_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  cin_IO_L2_in134_U0_fifo_cin_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    cin_IO_L2_in134_U0_fifo_cin_out_V_V_write_pass_0_q0 <= cin_IO_L2_in134_U0_fifo_cin_out_V_V_write_pass_0_out;
  end
  assign cin_IO_L2_in134_U0_fifo_cin_out_V_V_write_pass_0_in = cin_IO_L2_in134_U0_fifo_cin_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_5_9_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_5_9_V_V_full_n_pass_0_q0 <= fifo_w_PE_5_9_V_V_full_n_pass_0_out;
  end
  assign fifo_w_PE_5_9_V_V_full_n_pass_0_in = fifo_w_PE_5_9_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_cout_drain_IO_L1_out_9_5_V_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_cout_drain_IO_L1_out_9_5_V_V_full_n_pass_1_q0 <= fifo_cout_drain_cout_drain_IO_L1_out_9_5_V_V_full_n_pass_1_out;
  end
  assign fifo_cout_drain_cout_drain_IO_L1_out_9_5_V_V_full_n_pass_1_in = fifo_cout_drain_cout_drain_IO_L1_out_9_5_V_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg [31:0] PE_wrapper219_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper219_U0_fifo_cout_drain_out_V_din_pass_0_q0 <= PE_wrapper219_U0_fifo_cout_drain_out_V_din_pass_0_out;
  end
  assign PE_wrapper219_U0_fifo_cout_drain_out_V_din_pass_0_in = PE_wrapper219_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper219_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper219_U0_fifo_cout_drain_out_V_write_pass_0_q0 <= PE_wrapper219_U0_fifo_cout_drain_out_V_write_pass_0_out;
  end
  assign PE_wrapper219_U0_fifo_cout_drain_out_V_write_pass_0_in = PE_wrapper219_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  ap_done_Boundary_X6Y12_To_X8Y12_q0;
  always @ (posedge ap_clk) begin
    ap_done_Boundary_X6Y12_To_X8Y12_q0 <= ap_done_Boundary_X6Y12_To_X8Y12_out;
  end
  assign ap_done_Boundary_X6Y12_To_X8Y12_in = ap_done_Boundary_X6Y12_To_X8Y12_q0;
  (* dont_touch = "yes" *) reg  ap_start_Boundary_X6Y14_To_X8Y14_q0;
  always @ (posedge ap_clk) begin
    ap_start_Boundary_X6Y14_To_X8Y14_q0 <= ap_start_Boundary_X6Y14_To_X8Y14_out;
  end
  assign ap_start_Boundary_X6Y14_To_X8Y14_in = ap_start_Boundary_X6Y14_To_X8Y14_q0;
  (* dont_touch = "yes" *) reg  ap_rst_n_Boundary_X6Y14_To_X8Y14_q0;
  always @ (posedge ap_clk) begin
    ap_rst_n_Boundary_X6Y14_To_X8Y14_q0 <= ap_rst_n_Boundary_X6Y14_To_X8Y14_out;
  end
  assign ap_rst_n_Boundary_X6Y14_To_X8Y14_in = ap_rst_n_Boundary_X6Y14_To_X8Y14_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper231_U0_fifo_cin_out_V_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper231_U0_fifo_cin_out_V_V_din_pass_1_q0 <= PE_wrapper231_U0_fifo_cin_out_V_V_din_pass_1_out;
  end
  assign PE_wrapper231_U0_fifo_cin_out_V_V_din_pass_1_in = PE_wrapper231_U0_fifo_cin_out_V_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_7_9_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_7_9_V_V_full_n_pass_0_q0 <= fifo_cin_PE_7_9_V_V_full_n_pass_0_out;
  end
  assign fifo_cin_PE_7_9_V_V_full_n_pass_0_in = fifo_cin_PE_7_9_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper231_U0_fifo_cin_out_V_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper231_U0_fifo_cin_out_V_V_write_pass_1_q0 <= PE_wrapper231_U0_fifo_cin_out_V_V_write_pass_1_out;
  end
  assign PE_wrapper231_U0_fifo_cin_out_V_V_write_pass_1_in = PE_wrapper231_U0_fifo_cin_out_V_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [63:0] cout_drain_IO_L1_out_wrapper523_U0_fifo_cout_drain_out_V_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper523_U0_fifo_cout_drain_out_V_V_din_pass_1_q0 <= cout_drain_IO_L1_out_wrapper523_U0_fifo_cout_drain_out_V_V_din_pass_1_out;
  end
  assign cout_drain_IO_L1_out_wrapper523_U0_fifo_cout_drain_out_V_V_din_pass_1_in = cout_drain_IO_L1_out_wrapper523_U0_fifo_cout_drain_out_V_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_cout_drain_IO_L1_out_9_3_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_cout_drain_IO_L1_out_9_3_V_V_full_n_pass_0_q0 <= fifo_cout_drain_cout_drain_IO_L1_out_9_3_V_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_cout_drain_IO_L1_out_9_3_V_V_full_n_pass_0_in = fifo_cout_drain_cout_drain_IO_L1_out_9_3_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  cout_drain_IO_L1_out_wrapper523_U0_fifo_cout_drain_out_V_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper523_U0_fifo_cout_drain_out_V_V_write_pass_1_q0 <= cout_drain_IO_L1_out_wrapper523_U0_fifo_cout_drain_out_V_V_write_pass_1_out;
  end
  assign cout_drain_IO_L1_out_wrapper523_U0_fifo_cout_drain_out_V_V_write_pass_1_in = cout_drain_IO_L1_out_wrapper523_U0_fifo_cout_drain_out_V_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [63:0] cout_drain_IO_L2_out558_U0_fifo_cout_drain_out_V_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L2_out558_U0_fifo_cout_drain_out_V_V_din_pass_1_q0 <= cout_drain_IO_L2_out558_U0_fifo_cout_drain_out_V_V_din_pass_1_out;
  end
  assign cout_drain_IO_L2_out558_U0_fifo_cout_drain_out_V_V_din_pass_1_in = cout_drain_IO_L2_out558_U0_fifo_cout_drain_out_V_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_cout_drain_IO_L2_out_10_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_cout_drain_IO_L2_out_10_V_V_full_n_pass_0_q0 <= fifo_cout_drain_cout_drain_IO_L2_out_10_V_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_cout_drain_IO_L2_out_10_V_V_full_n_pass_0_in = fifo_cout_drain_cout_drain_IO_L2_out_10_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  cout_drain_IO_L2_out558_U0_fifo_cout_drain_out_V_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L2_out558_U0_fifo_cout_drain_out_V_V_write_pass_1_q0 <= cout_drain_IO_L2_out558_U0_fifo_cout_drain_out_V_V_write_pass_1_out;
  end
  assign cout_drain_IO_L2_out558_U0_fifo_cout_drain_out_V_V_write_pass_1_in = cout_drain_IO_L2_out558_U0_fifo_cout_drain_out_V_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper195_U0_fifo_cin_out_V_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper195_U0_fifo_cin_out_V_V_din_pass_1_q0 <= PE_wrapper195_U0_fifo_cin_out_V_V_din_pass_1_out;
  end
  assign PE_wrapper195_U0_fifo_cin_out_V_V_din_pass_1_in = PE_wrapper195_U0_fifo_cin_out_V_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_4_9_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_4_9_V_V_full_n_pass_0_q0 <= fifo_cin_PE_4_9_V_V_full_n_pass_0_out;
  end
  assign fifo_cin_PE_4_9_V_V_full_n_pass_0_in = fifo_cin_PE_4_9_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper195_U0_fifo_cin_out_V_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper195_U0_fifo_cin_out_V_V_write_pass_1_q0 <= PE_wrapper195_U0_fifo_cin_out_V_V_write_pass_1_out;
  end
  assign PE_wrapper195_U0_fifo_cin_out_V_V_write_pass_1_in = PE_wrapper195_U0_fifo_cin_out_V_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [63:0] cout_drain_IO_L1_out_wrapper521_U0_fifo_cout_drain_out_V_V_din_pass_1_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper521_U0_fifo_cout_drain_out_V_V_din_pass_1_q0 <= cout_drain_IO_L1_out_wrapper521_U0_fifo_cout_drain_out_V_V_din_pass_1_out;
  end
  assign cout_drain_IO_L1_out_wrapper521_U0_fifo_cout_drain_out_V_V_din_pass_1_in = cout_drain_IO_L1_out_wrapper521_U0_fifo_cout_drain_out_V_V_din_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_cout_drain_IO_L1_out_9_5_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_cout_drain_IO_L1_out_9_5_V_V_full_n_pass_0_q0 <= fifo_cout_drain_cout_drain_IO_L1_out_9_5_V_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_cout_drain_IO_L1_out_9_5_V_V_full_n_pass_0_in = fifo_cout_drain_cout_drain_IO_L1_out_9_5_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  cout_drain_IO_L1_out_wrapper521_U0_fifo_cout_drain_out_V_V_write_pass_1_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper521_U0_fifo_cout_drain_out_V_V_write_pass_1_q0 <= cout_drain_IO_L1_out_wrapper521_U0_fifo_cout_drain_out_V_V_write_pass_1_out;
  end
  assign cout_drain_IO_L1_out_wrapper521_U0_fifo_cout_drain_out_V_V_write_pass_1_in = cout_drain_IO_L1_out_wrapper521_U0_fifo_cout_drain_out_V_V_write_pass_1_q0;
  (* dont_touch = "yes" *) reg [63:0] cout_drain_IO_L1_out_wrapper551_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper551_U0_fifo_cout_drain_out_V_V_din_pass_0_q0 <= cout_drain_IO_L1_out_wrapper551_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper551_U0_fifo_cout_drain_out_V_V_din_pass_0_in = cout_drain_IO_L1_out_wrapper551_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  cout_drain_IO_L1_out_wrapper551_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper551_U0_fifo_cout_drain_out_V_V_write_pass_0_q0 <= cout_drain_IO_L1_out_wrapper551_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper551_U0_fifo_cout_drain_out_V_V_write_pass_0_in = cout_drain_IO_L1_out_wrapper551_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_cout_drain_IO_L1_out_11_1_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_cout_drain_IO_L1_out_11_1_V_V_full_n_pass_0_q0 <= fifo_cout_drain_cout_drain_IO_L1_out_11_1_V_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_cout_drain_IO_L1_out_11_1_V_V_full_n_pass_0_in = fifo_cout_drain_cout_drain_IO_L1_out_11_1_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_0_11_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_0_11_V_V_full_n_pass_0_q0 <= fifo_w_PE_0_11_V_V_full_n_pass_0_out;
  end
  assign fifo_w_PE_0_11_V_V_full_n_pass_0_in = fifo_w_PE_0_11_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_8_10_V_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_8_10_V_V_full_n_pass_1_q0 <= fifo_cin_PE_8_10_V_V_full_n_pass_1_out;
  end
  assign fifo_cin_PE_8_10_V_V_full_n_pass_1_in = fifo_cin_PE_8_10_V_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_1_12_V_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_1_12_V_V_full_n_pass_1_q0 <= fifo_w_PE_1_12_V_V_full_n_pass_1_out;
  end
  assign fifo_w_PE_1_12_V_V_full_n_pass_1_in = fifo_w_PE_1_12_V_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_2_11_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_2_11_V_V_full_n_pass_0_q0 <= fifo_w_PE_2_11_V_V_full_n_pass_0_out;
  end
  assign fifo_w_PE_2_11_V_V_full_n_pass_0_in = fifo_w_PE_2_11_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper161_U0_fifo_cin_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper161_U0_fifo_cin_out_V_V_din_pass_0_q0 <= PE_wrapper161_U0_fifo_cin_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper161_U0_fifo_cin_out_V_V_din_pass_0_in = PE_wrapper161_U0_fifo_cin_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper161_U0_fifo_cin_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper161_U0_fifo_cin_out_V_V_write_pass_0_q0 <= PE_wrapper161_U0_fifo_cin_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper161_U0_fifo_cin_out_V_V_write_pass_0_in = PE_wrapper161_U0_fifo_cin_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper256_U0_fifo_cin_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper256_U0_fifo_cin_out_V_V_din_pass_0_q0 <= PE_wrapper256_U0_fifo_cin_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper256_U0_fifo_cin_out_V_V_din_pass_0_in = PE_wrapper256_U0_fifo_cin_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper256_U0_fifo_cin_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper256_U0_fifo_cin_out_V_V_write_pass_0_q0 <= PE_wrapper256_U0_fifo_cin_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper256_U0_fifo_cin_out_V_V_write_pass_0_in = PE_wrapper256_U0_fifo_cin_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_3_11_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_3_11_V_V_full_n_pass_0_q0 <= fifo_w_PE_3_11_V_V_full_n_pass_0_out;
  end
  assign fifo_w_PE_3_11_V_V_full_n_pass_0_in = fifo_w_PE_3_11_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_4_12_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_4_12_V_V_full_n_pass_0_q0 <= fifo_w_PE_4_12_V_V_full_n_pass_0_out;
  end
  assign fifo_w_PE_4_12_V_V_full_n_pass_0_in = fifo_w_PE_4_12_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_7_11_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_7_11_V_V_full_n_pass_0_q0 <= fifo_cin_PE_7_11_V_V_full_n_pass_0_out;
  end
  assign fifo_cin_PE_7_11_V_V_full_n_pass_0_in = fifo_cin_PE_7_11_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_PE_8_9_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_PE_8_9_V_full_n_pass_1_q0 <= fifo_cout_drain_PE_8_9_V_full_n_pass_1_out;
  end
  assign fifo_cout_drain_PE_8_9_V_full_n_pass_1_in = fifo_cout_drain_PE_8_9_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper197_U0_fifo_cin_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper197_U0_fifo_cin_out_V_V_din_pass_0_q0 <= PE_wrapper197_U0_fifo_cin_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper197_U0_fifo_cin_out_V_V_din_pass_0_in = PE_wrapper197_U0_fifo_cin_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper197_U0_fifo_cin_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper197_U0_fifo_cin_out_V_V_write_pass_0_q0 <= PE_wrapper197_U0_fifo_cin_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper197_U0_fifo_cin_out_V_V_write_pass_0_in = PE_wrapper197_U0_fifo_cin_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [31:0] PE_wrapper185_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper185_U0_fifo_cout_drain_out_V_din_pass_0_q0 <= PE_wrapper185_U0_fifo_cout_drain_out_V_din_pass_0_out;
  end
  assign PE_wrapper185_U0_fifo_cout_drain_out_V_din_pass_0_in = PE_wrapper185_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper185_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper185_U0_fifo_cout_drain_out_V_write_pass_0_q0 <= PE_wrapper185_U0_fifo_cout_drain_out_V_write_pass_0_out;
  end
  assign PE_wrapper185_U0_fifo_cout_drain_out_V_write_pass_0_in = PE_wrapper185_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [63:0] cout_drain_IO_L1_out_wrapper518_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper518_U0_fifo_cout_drain_out_V_V_din_pass_0_q0 <= cout_drain_IO_L1_out_wrapper518_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper518_U0_fifo_cout_drain_out_V_V_din_pass_0_in = cout_drain_IO_L1_out_wrapper518_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  cout_drain_IO_L1_out_wrapper518_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper518_U0_fifo_cout_drain_out_V_V_write_pass_0_q0 <= cout_drain_IO_L1_out_wrapper518_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper518_U0_fifo_cout_drain_out_V_V_write_pass_0_in = cout_drain_IO_L1_out_wrapper518_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_7_11_V_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_7_11_V_V_full_n_pass_1_q0 <= fifo_w_PE_7_11_V_V_full_n_pass_1_out;
  end
  assign fifo_w_PE_7_11_V_V_full_n_pass_1_in = fifo_w_PE_7_11_V_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_cout_drain_IO_L1_out_9_9_V_V_full_n_pass_2_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_cout_drain_IO_L1_out_9_9_V_V_full_n_pass_2_q0 <= fifo_cout_drain_cout_drain_IO_L1_out_9_9_V_V_full_n_pass_2_out;
  end
  assign fifo_cout_drain_cout_drain_IO_L1_out_9_9_V_V_full_n_pass_2_in = fifo_cout_drain_cout_drain_IO_L1_out_9_9_V_V_full_n_pass_2_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_cout_drain_IO_L1_out_11_8_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_cout_drain_IO_L1_out_11_8_V_V_full_n_pass_0_q0 <= fifo_cout_drain_cout_drain_IO_L1_out_11_8_V_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_cout_drain_IO_L1_out_11_8_V_V_full_n_pass_0_in = fifo_cout_drain_cout_drain_IO_L1_out_11_8_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_w_PE_8_10_V_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_w_PE_8_10_V_V_full_n_pass_1_q0 <= fifo_w_PE_8_10_V_V_full_n_pass_1_out;
  end
  assign fifo_w_PE_8_10_V_V_full_n_pass_1_in = fifo_w_PE_8_10_V_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg [63:0] cout_drain_IO_L1_out_wrapper534_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper534_U0_fifo_cout_drain_out_V_V_din_pass_0_q0 <= cout_drain_IO_L1_out_wrapper534_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper534_U0_fifo_cout_drain_out_V_V_din_pass_0_in = cout_drain_IO_L1_out_wrapper534_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  cout_drain_IO_L1_out_wrapper534_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L1_out_wrapper534_U0_fifo_cout_drain_out_V_V_write_pass_0_q0 <= cout_drain_IO_L1_out_wrapper534_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  end
  assign cout_drain_IO_L1_out_wrapper534_U0_fifo_cout_drain_out_V_V_write_pass_0_in = cout_drain_IO_L1_out_wrapper534_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper257_U0_fifo_cin_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper257_U0_fifo_cin_out_V_V_din_pass_0_q0 <= PE_wrapper257_U0_fifo_cin_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper257_U0_fifo_cin_out_V_V_din_pass_0_in = PE_wrapper257_U0_fifo_cin_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper257_U0_fifo_cin_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper257_U0_fifo_cin_out_V_V_write_pass_0_q0 <= PE_wrapper257_U0_fifo_cin_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper257_U0_fifo_cin_out_V_V_write_pass_0_in = PE_wrapper257_U0_fifo_cin_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [31:0] PE_wrapper257_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper257_U0_fifo_cout_drain_out_V_din_pass_0_q0 <= PE_wrapper257_U0_fifo_cout_drain_out_V_din_pass_0_out;
  end
  assign PE_wrapper257_U0_fifo_cout_drain_out_V_din_pass_0_in = PE_wrapper257_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper257_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper257_U0_fifo_cout_drain_out_V_write_pass_0_q0 <= PE_wrapper257_U0_fifo_cout_drain_out_V_write_pass_0_out;
  end
  assign PE_wrapper257_U0_fifo_cout_drain_out_V_write_pass_0_in = PE_wrapper257_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_0_11_V_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_0_11_V_V_full_n_pass_0_q0 <= fifo_cin_PE_0_11_V_V_full_n_pass_0_out;
  end
  assign fifo_cin_PE_0_11_V_V_full_n_pass_0_in = fifo_cin_PE_0_11_V_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cin_PE_2_11_V_V_full_n_pass_1_q0;
  always @ (posedge ap_clk) begin
    fifo_cin_PE_2_11_V_V_full_n_pass_1_q0 <= fifo_cin_PE_2_11_V_V_full_n_pass_1_out;
  end
  assign fifo_cin_PE_2_11_V_V_full_n_pass_1_in = fifo_cin_PE_2_11_V_V_full_n_pass_1_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_cout_drain_IO_L1_out_10_9_V_V_full_n_pass_2_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_cout_drain_IO_L1_out_10_9_V_V_full_n_pass_2_q0 <= fifo_cout_drain_cout_drain_IO_L1_out_10_9_V_V_full_n_pass_2_out;
  end
  assign fifo_cout_drain_cout_drain_IO_L1_out_10_9_V_V_full_n_pass_2_in = fifo_cout_drain_cout_drain_IO_L1_out_10_9_V_V_full_n_pass_2_q0;
  (* dont_touch = "yes" *) reg [31:0] PE_wrapper197_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper197_U0_fifo_cout_drain_out_V_din_pass_0_q0 <= PE_wrapper197_U0_fifo_cout_drain_out_V_din_pass_0_out;
  end
  assign PE_wrapper197_U0_fifo_cout_drain_out_V_din_pass_0_in = PE_wrapper197_U0_fifo_cout_drain_out_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper197_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper197_U0_fifo_cout_drain_out_V_write_pass_0_q0 <= PE_wrapper197_U0_fifo_cout_drain_out_V_write_pass_0_out;
  end
  assign PE_wrapper197_U0_fifo_cout_drain_out_V_write_pass_0_in = PE_wrapper197_U0_fifo_cout_drain_out_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  fifo_cout_drain_PE_6_11_V_full_n_pass_0_q0;
  always @ (posedge ap_clk) begin
    fifo_cout_drain_PE_6_11_V_full_n_pass_0_q0 <= fifo_cout_drain_PE_6_11_V_full_n_pass_0_out;
  end
  assign fifo_cout_drain_PE_6_11_V_full_n_pass_0_in = fifo_cout_drain_PE_6_11_V_full_n_pass_0_q0;
  (* dont_touch = "yes" *) reg [255:0] PE_wrapper185_U0_fifo_w_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper185_U0_fifo_w_out_V_V_din_pass_0_q0 <= PE_wrapper185_U0_fifo_w_out_V_V_din_pass_0_out;
  end
  assign PE_wrapper185_U0_fifo_w_out_V_V_din_pass_0_in = PE_wrapper185_U0_fifo_w_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  PE_wrapper185_U0_fifo_w_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    PE_wrapper185_U0_fifo_w_out_V_V_write_pass_0_q0 <= PE_wrapper185_U0_fifo_w_out_V_V_write_pass_0_out;
  end
  assign PE_wrapper185_U0_fifo_w_out_V_V_write_pass_0_in = PE_wrapper185_U0_fifo_w_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg [63:0] cout_drain_IO_L2_out_boundary_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L2_out_boundary_U0_fifo_cout_drain_out_V_V_din_pass_0_q0 <= cout_drain_IO_L2_out_boundary_U0_fifo_cout_drain_out_V_V_din_pass_0_out;
  end
  assign cout_drain_IO_L2_out_boundary_U0_fifo_cout_drain_out_V_V_din_pass_0_in = cout_drain_IO_L2_out_boundary_U0_fifo_cout_drain_out_V_V_din_pass_0_q0;
  (* dont_touch = "yes" *) reg  cout_drain_IO_L2_out_boundary_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  always @ (posedge ap_clk) begin
    cout_drain_IO_L2_out_boundary_U0_fifo_cout_drain_out_V_V_write_pass_0_q0 <= cout_drain_IO_L2_out_boundary_U0_fifo_cout_drain_out_V_V_write_pass_0_out;
  end
  assign cout_drain_IO_L2_out_boundary_U0_fifo_cout_drain_out_V_V_write_pass_0_in = cout_drain_IO_L2_out_boundary_U0_fifo_cout_drain_out_V_V_write_pass_0_q0;
  (* dont_touch = "yes" *) reg  ap_done_Boundary_X6Y14_To_X8Y14_q0;
  always @ (posedge ap_clk) begin
    ap_done_Boundary_X6Y14_To_X8Y14_q0 <= ap_done_Boundary_X6Y14_To_X8Y14_out;
  end
  assign ap_done_Boundary_X6Y14_To_X8Y14_in = ap_done_Boundary_X6Y14_To_X8Y14_q0;
wire ap_done = ap_done_Boundary_X4Y2_To_X6Y2_in & ap_done_Boundary_X6Y0_To_X6Y2_in & ap_done_Boundary_X4Y0_To_X4Y2_in;
wire ap_idle = ap_done;
wire ap_ready = ap_done;
wire ap_start = ap_start_Boundary_X4Y2_To_X6Y2_out;


  (* keep_hierarchy = "yes" *) CR_X4Y0_To_CR_X5Y1_ctrl CR_X4Y0_To_CR_X5Y1_ctrl_U0 (
    .PE_wrapper211_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper211_U0_fifo_cin_out_V_V_din_pass_0_in),
    .PE_wrapper211_U0_fifo_cin_out_V_V_din_pass_1(PE_wrapper211_U0_fifo_cin_out_V_V_din_pass_1_out),
    .fifo_cin_PE_6_1_V_V_full_n_pass_0(fifo_cin_PE_6_1_V_V_full_n_pass_0_out),
    .fifo_cin_PE_6_1_V_V_full_n_pass_1(fifo_cin_PE_6_1_V_V_full_n_pass_1_in),
    .PE_wrapper211_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper211_U0_fifo_cin_out_V_V_write_pass_0_in),
    .PE_wrapper211_U0_fifo_cin_out_V_V_write_pass_1(PE_wrapper211_U0_fifo_cin_out_V_V_write_pass_1_out),
    .PE_wrapper212_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper212_U0_fifo_cin_out_V_V_din_pass_0_in),
    .PE_wrapper212_U0_fifo_cin_out_V_V_din_pass_1(PE_wrapper212_U0_fifo_cin_out_V_V_din_pass_1_out),
    .fifo_cin_PE_6_2_V_V_full_n_pass_0(fifo_cin_PE_6_2_V_V_full_n_pass_0_out),
    .fifo_cin_PE_6_2_V_V_full_n_pass_1(fifo_cin_PE_6_2_V_V_full_n_pass_1_in),
    .PE_wrapper212_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper212_U0_fifo_cin_out_V_V_write_pass_0_in),
    .PE_wrapper212_U0_fifo_cin_out_V_V_write_pass_1(PE_wrapper212_U0_fifo_cin_out_V_V_write_pass_1_out),
    .PE_wrapper213_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper213_U0_fifo_cin_out_V_V_din_pass_0_in),
    .PE_wrapper213_U0_fifo_cin_out_V_V_din_pass_1(PE_wrapper213_U0_fifo_cin_out_V_V_din_pass_1_out),
    .fifo_cin_PE_6_3_V_V_full_n_pass_0(fifo_cin_PE_6_3_V_V_full_n_pass_0_out),
    .fifo_cin_PE_6_3_V_V_full_n_pass_1(fifo_cin_PE_6_3_V_V_full_n_pass_1_in),
    .PE_wrapper213_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper213_U0_fifo_cin_out_V_V_write_pass_0_in),
    .PE_wrapper213_U0_fifo_cin_out_V_V_write_pass_1(PE_wrapper213_U0_fifo_cin_out_V_V_write_pass_1_out),
    .cin_IO_L2_in125_U0_fifo_cin_out_V_V_din_pass_0(cin_IO_L2_in125_U0_fifo_cin_out_V_V_din_pass_0_in),
    .cin_IO_L2_in125_U0_fifo_cin_out_V_V_din_pass_1(cin_IO_L2_in125_U0_fifo_cin_out_V_V_din_pass_1_out),
    .fifo_cin_cin_IO_L2_in_2_V_V_full_n_pass_0(fifo_cin_cin_IO_L2_in_2_V_V_full_n_pass_0_out),
    .fifo_cin_cin_IO_L2_in_2_V_V_full_n_pass_1(fifo_cin_cin_IO_L2_in_2_V_V_full_n_pass_1_in),
    .cin_IO_L2_in125_U0_fifo_cin_out_V_V_write_pass_0(cin_IO_L2_in125_U0_fifo_cin_out_V_V_write_pass_0_in),
    .cin_IO_L2_in125_U0_fifo_cin_out_V_V_write_pass_1(cin_IO_L2_in125_U0_fifo_cin_out_V_V_write_pass_1_out),
    .cout_drain_IO_L1_out_wrapper424_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper424_U0_fifo_cout_drain_out_V_V_din_pass_0_in),
    .cout_drain_IO_L1_out_wrapper424_U0_fifo_cout_drain_out_V_V_din_pass_1(cout_drain_IO_L1_out_wrapper424_U0_fifo_cout_drain_out_V_V_din_pass_1_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_3_6_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_3_6_V_V_full_n_pass_0_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_3_6_V_V_full_n_pass_1(fifo_cout_drain_cout_drain_IO_L1_out_3_6_V_V_full_n_pass_1_in),
    .cout_drain_IO_L1_out_wrapper424_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper424_U0_fifo_cout_drain_out_V_V_write_pass_0_in),
    .cout_drain_IO_L1_out_wrapper424_U0_fifo_cout_drain_out_V_V_write_pass_1(cout_drain_IO_L1_out_wrapper424_U0_fifo_cout_drain_out_V_V_write_pass_1_out),
    .cout_drain_IO_L1_out_wrapper408_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper408_U0_fifo_cout_drain_out_V_V_din_pass_0_in),
    .cout_drain_IO_L1_out_wrapper408_U0_fifo_cout_drain_out_V_V_din_pass_1(cout_drain_IO_L1_out_wrapper408_U0_fifo_cout_drain_out_V_V_din_pass_1_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_2_6_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_2_6_V_V_full_n_pass_0_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_2_6_V_V_full_n_pass_1(fifo_cout_drain_cout_drain_IO_L1_out_2_6_V_V_full_n_pass_1_in),
    .cout_drain_IO_L1_out_wrapper408_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper408_U0_fifo_cout_drain_out_V_V_write_pass_0_in),
    .cout_drain_IO_L1_out_wrapper408_U0_fifo_cout_drain_out_V_V_write_pass_1(cout_drain_IO_L1_out_wrapper408_U0_fifo_cout_drain_out_V_V_write_pass_1_out),
    .cout_drain_IO_L1_out_wrapper376_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper376_U0_fifo_cout_drain_out_V_V_din_pass_0_in),
    .cout_drain_IO_L1_out_wrapper376_U0_fifo_cout_drain_out_V_V_din_pass_1(cout_drain_IO_L1_out_wrapper376_U0_fifo_cout_drain_out_V_V_din_pass_1_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_0_6_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_0_6_V_V_full_n_pass_0_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_0_6_V_V_full_n_pass_1(fifo_cout_drain_cout_drain_IO_L1_out_0_6_V_V_full_n_pass_1_in),
    .cout_drain_IO_L1_out_wrapper376_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper376_U0_fifo_cout_drain_out_V_V_write_pass_0_in),
    .cout_drain_IO_L1_out_wrapper376_U0_fifo_cout_drain_out_V_V_write_pass_1(cout_drain_IO_L1_out_wrapper376_U0_fifo_cout_drain_out_V_V_write_pass_1_out),
    .cout_drain_IO_L1_out_wrapper392_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper392_U0_fifo_cout_drain_out_V_V_din_pass_0_in),
    .cout_drain_IO_L1_out_wrapper392_U0_fifo_cout_drain_out_V_V_din_pass_1(cout_drain_IO_L1_out_wrapper392_U0_fifo_cout_drain_out_V_V_din_pass_1_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_1_6_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_1_6_V_V_full_n_pass_0_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_1_6_V_V_full_n_pass_1(fifo_cout_drain_cout_drain_IO_L1_out_1_6_V_V_full_n_pass_1_in),
    .cout_drain_IO_L1_out_wrapper392_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper392_U0_fifo_cout_drain_out_V_V_write_pass_0_in),
    .cout_drain_IO_L1_out_wrapper392_U0_fifo_cout_drain_out_V_V_write_pass_1(cout_drain_IO_L1_out_wrapper392_U0_fifo_cout_drain_out_V_V_write_pass_1_out),
    .PE_wrapper213_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper213_U0_fifo_w_out_V_V_din_pass_0_in),
    .PE_wrapper213_U0_fifo_w_out_V_V_din_pass_1(PE_wrapper213_U0_fifo_w_out_V_V_din_pass_1_out),
    .fifo_w_PE_5_4_V_V_full_n_pass_0(fifo_w_PE_5_4_V_V_full_n_pass_0_out),
    .fifo_w_PE_5_4_V_V_full_n_pass_1(fifo_w_PE_5_4_V_V_full_n_pass_1_in),
    .PE_wrapper213_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper213_U0_fifo_w_out_V_V_write_pass_0_in),
    .PE_wrapper213_U0_fifo_w_out_V_V_write_pass_1(PE_wrapper213_U0_fifo_w_out_V_V_write_pass_1_out),
    .PE_wrapper187_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper187_U0_fifo_w_out_V_V_din_pass_0_out),
    .fifo_w_PE_3_2_V_V_full_n_pass_0(fifo_w_PE_3_2_V_V_full_n_pass_0_in),
    .PE_wrapper187_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper187_U0_fifo_w_out_V_V_write_pass_0_out),
    .PE_wrapper187_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper187_U0_fifo_cout_drain_out_V_din_pass_0_out),
    .fifo_cout_drain_PE_3_1_V_full_n_pass_0(fifo_cout_drain_PE_3_1_V_full_n_pass_0_in),
    .PE_wrapper187_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper187_U0_fifo_cout_drain_out_V_write_pass_0_out),
    .PE_wrapper162_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper162_U0_fifo_cin_out_V_V_din_pass_0_in),
    .fifo_cin_PE_2_0_V_V_full_n_pass_0(fifo_cin_PE_2_0_V_V_full_n_pass_0_out),
    .PE_wrapper162_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper162_U0_fifo_cin_out_V_V_write_pass_0_in),
    .w_IO_L2_in137_U0_fifo_w_out_V_V_din_pass_0(w_IO_L2_in137_U0_fifo_w_out_V_V_din_pass_0_out),
    .fifo_w_w_IO_L2_in_3_V_V_full_n_pass_0(fifo_w_w_IO_L2_in_3_V_V_full_n_pass_0_in),
    .w_IO_L2_in137_U0_fifo_w_out_V_V_write_pass_0(w_IO_L2_in137_U0_fifo_w_out_V_V_write_pass_0_out),
    .PE_wrapper151_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper151_U0_fifo_cout_drain_out_V_din_pass_0_out),
    .fifo_cout_drain_PE_0_1_V_full_n_pass_0(fifo_cout_drain_PE_0_1_V_full_n_pass_0_in),
    .PE_wrapper151_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper151_U0_fifo_cout_drain_out_V_write_pass_0_out),
    .PE_wrapper163_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper163_U0_fifo_w_out_V_V_din_pass_0_out),
    .fifo_w_PE_1_2_V_V_full_n_pass_0(fifo_w_PE_1_2_V_V_full_n_pass_0_in),
    .PE_wrapper163_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper163_U0_fifo_w_out_V_V_write_pass_0_out),
    .w_IO_L2_in136_U0_fifo_w_out_V_V_din_pass_0(w_IO_L2_in136_U0_fifo_w_out_V_V_din_pass_0_in),
    .fifo_w_w_IO_L2_in_2_V_V_full_n_pass_0(fifo_w_w_IO_L2_in_2_V_V_full_n_pass_0_out),
    .w_IO_L2_in136_U0_fifo_w_out_V_V_write_pass_0(w_IO_L2_in136_U0_fifo_w_out_V_V_write_pass_0_in),
    .cin_IO_L2_in124_U0_fifo_cin_out_V_V_din_pass_0(cin_IO_L2_in124_U0_fifo_cin_out_V_V_din_pass_0_out),
    .fifo_cin_cin_IO_L2_in_1_V_V_full_n_pass_0(fifo_cin_cin_IO_L2_in_1_V_V_full_n_pass_0_in),
    .cin_IO_L2_in124_U0_fifo_cin_out_V_V_write_pass_0(cin_IO_L2_in124_U0_fifo_cin_out_V_V_write_pass_0_out),
    .w_IO_L2_in138_U0_fifo_w_local_out_V_V_din_pass_1(w_IO_L2_in138_U0_fifo_w_local_out_V_V_din_pass_1_in),
    .fifo_w_PE_3_0_V_V_full_n_pass_1(fifo_w_PE_3_0_V_V_full_n_pass_1_out),
    .w_IO_L2_in138_U0_fifo_w_local_out_V_V_write_pass_1(w_IO_L2_in138_U0_fifo_w_local_out_V_V_write_pass_1_in),
    .kernel0_entry12_U0_w_V_out_din_pass_0(kernel0_entry12_U0_w_V_out_din_pass_0_out),
    .w_V_c_full_n_pass_0(w_V_c_full_n_pass_0_in),
    .kernel0_entry12_U0_w_V_out_write_pass_0(kernel0_entry12_U0_w_V_out_write_pass_0_out),
    .PE_wrapper163_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper163_U0_fifo_cout_drain_out_V_din_pass_0_out),
    .fifo_cout_drain_PE_1_1_V_full_n_pass_0(fifo_cout_drain_PE_1_1_V_full_n_pass_0_in),
    .PE_wrapper163_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper163_U0_fifo_cout_drain_out_V_write_pass_0_out),
    .PE_wrapper151_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper151_U0_fifo_w_out_V_V_din_pass_0_out),
    .fifo_w_PE_0_2_V_V_full_n_pass_0(fifo_w_PE_0_2_V_V_full_n_pass_0_in),
    .PE_wrapper151_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper151_U0_fifo_w_out_V_V_write_pass_0_out),
    .PE_wrapper162_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper162_U0_fifo_cout_drain_out_V_din_pass_0_in),
    .fifo_cout_drain_PE_1_0_V_full_n_pass_0(fifo_cout_drain_PE_1_0_V_full_n_pass_0_out),
    .PE_wrapper162_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper162_U0_fifo_cout_drain_out_V_write_pass_0_in),
    .PE_wrapper150_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper150_U0_fifo_cin_out_V_V_din_pass_0_out),
    .fifo_cin_PE_1_0_V_V_full_n_pass_0(fifo_cin_PE_1_0_V_V_full_n_pass_0_in),
    .PE_wrapper150_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper150_U0_fifo_cin_out_V_V_write_pass_0_out),
    .PE_wrapper175_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper175_U0_fifo_cout_drain_out_V_din_pass_0_out),
    .fifo_cout_drain_PE_2_1_V_full_n_pass_0(fifo_cout_drain_PE_2_1_V_full_n_pass_0_in),
    .PE_wrapper175_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper175_U0_fifo_cout_drain_out_V_write_pass_0_out),
    .PE_wrapper175_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper175_U0_fifo_w_out_V_V_din_pass_0_out),
    .fifo_w_PE_2_2_V_V_full_n_pass_0(fifo_w_PE_2_2_V_V_full_n_pass_0_in),
    .PE_wrapper175_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper175_U0_fifo_w_out_V_V_write_pass_0_out),
    .cin_IO_L2_in125_U0_fifo_cin_local_out_V_V_din_pass_0(cin_IO_L2_in125_U0_fifo_cin_local_out_V_V_din_pass_0_in),
    .fifo_cin_PE_0_1_V_V_full_n_pass_0(fifo_cin_PE_0_1_V_V_full_n_pass_0_out),
    .cin_IO_L2_in125_U0_fifo_cin_local_out_V_V_write_pass_0(cin_IO_L2_in125_U0_fifo_cin_local_out_V_V_write_pass_0_in),
    .cout_drain_IO_L1_out_wrapper378_U0_fifo_cout_drain_out_V_V_din_pass_1(cout_drain_IO_L1_out_wrapper378_U0_fifo_cout_drain_out_V_V_din_pass_1_in),
    .fifo_cout_drain_cout_drain_IO_L1_out_0_4_V_V_full_n_pass_1(fifo_cout_drain_cout_drain_IO_L1_out_0_4_V_V_full_n_pass_1_out),
    .cout_drain_IO_L1_out_wrapper378_U0_fifo_cout_drain_out_V_V_write_pass_1(cout_drain_IO_L1_out_wrapper378_U0_fifo_cout_drain_out_V_V_write_pass_1_in),
    .kernel0_entry12_U0_cout_V_out_din_pass_0(kernel0_entry12_U0_cout_V_out_din_pass_0_out),
    .cout_V_c_full_n_pass_0(cout_V_c_full_n_pass_0_in),
    .kernel0_entry12_U0_cout_V_out_write_pass_0(kernel0_entry12_U0_cout_V_out_write_pass_0_out),
    .PE_wrapper187_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper187_U0_fifo_cin_out_V_V_din_pass_0_out),
    .fifo_cin_PE_4_1_V_V_full_n_pass_0(fifo_cin_PE_4_1_V_V_full_n_pass_0_in),
    .PE_wrapper187_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper187_U0_fifo_cin_out_V_V_write_pass_0_out),
    .PE_wrapper162_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper162_U0_fifo_w_out_V_V_din_pass_0_in),
    .fifo_w_PE_1_1_V_V_full_n_pass_0(fifo_w_PE_1_1_V_V_full_n_pass_0_out),
    .PE_wrapper162_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper162_U0_fifo_w_out_V_V_write_pass_0_in),
    .cout_drain_IO_L1_out_wrapper382_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper382_U0_fifo_cout_drain_out_V_V_din_pass_0_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_0_0_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_0_0_V_V_full_n_pass_0_in),
    .cout_drain_IO_L1_out_wrapper382_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper382_U0_fifo_cout_drain_out_V_V_write_pass_0_out),
    .PE_wrapper186_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper186_U0_fifo_cin_out_V_V_din_pass_0_out),
    .fifo_cin_PE_4_0_V_V_full_n_pass_0(fifo_cin_PE_4_0_V_V_full_n_pass_0_in),
    .PE_wrapper186_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper186_U0_fifo_cin_out_V_V_write_pass_0_out),
    .w_IO_L2_in135_U0_fifo_w_local_out_V_V_din_pass_0(w_IO_L2_in135_U0_fifo_w_local_out_V_V_din_pass_0_in),
    .fifo_w_PE_0_0_V_V_full_n_pass_0(fifo_w_PE_0_0_V_V_full_n_pass_0_out),
    .w_IO_L2_in135_U0_fifo_w_local_out_V_V_write_pass_0(w_IO_L2_in135_U0_fifo_w_local_out_V_V_write_pass_0_in),
    .s_axi_control_AWVALID(s_axi_control_AWVALID),
    .s_axi_control_AWREADY(s_axi_control_AWREADY),
    .s_axi_control_AWADDR(s_axi_control_AWADDR),
    .s_axi_control_WVALID(s_axi_control_WVALID),
    .s_axi_control_WREADY(s_axi_control_WREADY),
    .s_axi_control_WDATA(s_axi_control_WDATA),
    .s_axi_control_WSTRB(s_axi_control_WSTRB),
    .s_axi_control_ARVALID(s_axi_control_ARVALID),
    .s_axi_control_ARREADY(s_axi_control_ARREADY),
    .s_axi_control_ARADDR(s_axi_control_ARADDR),
    .s_axi_control_RVALID(s_axi_control_RVALID),
    .s_axi_control_RREADY(s_axi_control_RREADY),
    .s_axi_control_RDATA(s_axi_control_RDATA),
    .s_axi_control_RRESP(s_axi_control_RRESP),
    .s_axi_control_BVALID(s_axi_control_BVALID),
    .s_axi_control_BREADY(s_axi_control_BREADY),
    .s_axi_control_BRESP(s_axi_control_BRESP),
    .interrupt(interrupt),
    .m_axi_gmem_cin_AWVALID(m_axi_gmem_cin_AWVALID),
    .m_axi_gmem_cin_AWREADY(m_axi_gmem_cin_AWREADY),
    .m_axi_gmem_cin_AWADDR(m_axi_gmem_cin_AWADDR),
    .m_axi_gmem_cin_AWID(m_axi_gmem_cin_AWID),
    .m_axi_gmem_cin_AWLEN(m_axi_gmem_cin_AWLEN),
    .m_axi_gmem_cin_AWSIZE(m_axi_gmem_cin_AWSIZE),
    .m_axi_gmem_cin_AWBURST(m_axi_gmem_cin_AWBURST),
    .m_axi_gmem_cin_AWLOCK(m_axi_gmem_cin_AWLOCK),
    .m_axi_gmem_cin_AWCACHE(m_axi_gmem_cin_AWCACHE),
    .m_axi_gmem_cin_AWPROT(m_axi_gmem_cin_AWPROT),
    .m_axi_gmem_cin_AWQOS(m_axi_gmem_cin_AWQOS),
    .m_axi_gmem_cin_AWREGION(m_axi_gmem_cin_AWREGION),
    .m_axi_gmem_cin_AWUSER(m_axi_gmem_cin_AWUSER),
    .m_axi_gmem_cin_WVALID(m_axi_gmem_cin_WVALID),
    .m_axi_gmem_cin_WREADY(m_axi_gmem_cin_WREADY),
    .m_axi_gmem_cin_WDATA(m_axi_gmem_cin_WDATA),
    .m_axi_gmem_cin_WSTRB(m_axi_gmem_cin_WSTRB),
    .m_axi_gmem_cin_WLAST(m_axi_gmem_cin_WLAST),
    .m_axi_gmem_cin_WID(m_axi_gmem_cin_WID),
    .m_axi_gmem_cin_WUSER(m_axi_gmem_cin_WUSER),
    .m_axi_gmem_cin_ARVALID(m_axi_gmem_cin_ARVALID),
    .m_axi_gmem_cin_ARREADY(m_axi_gmem_cin_ARREADY),
    .m_axi_gmem_cin_ARADDR(m_axi_gmem_cin_ARADDR),
    .m_axi_gmem_cin_ARID(m_axi_gmem_cin_ARID),
    .m_axi_gmem_cin_ARLEN(m_axi_gmem_cin_ARLEN),
    .m_axi_gmem_cin_ARSIZE(m_axi_gmem_cin_ARSIZE),
    .m_axi_gmem_cin_ARBURST(m_axi_gmem_cin_ARBURST),
    .m_axi_gmem_cin_ARLOCK(m_axi_gmem_cin_ARLOCK),
    .m_axi_gmem_cin_ARCACHE(m_axi_gmem_cin_ARCACHE),
    .m_axi_gmem_cin_ARPROT(m_axi_gmem_cin_ARPROT),
    .m_axi_gmem_cin_ARQOS(m_axi_gmem_cin_ARQOS),
    .m_axi_gmem_cin_ARREGION(m_axi_gmem_cin_ARREGION),
    .m_axi_gmem_cin_ARUSER(m_axi_gmem_cin_ARUSER),
    .m_axi_gmem_cin_RVALID(m_axi_gmem_cin_RVALID),
    .m_axi_gmem_cin_RREADY(m_axi_gmem_cin_RREADY),
    .m_axi_gmem_cin_RDATA(m_axi_gmem_cin_RDATA),
    .m_axi_gmem_cin_RLAST(m_axi_gmem_cin_RLAST),
    .m_axi_gmem_cin_RID(m_axi_gmem_cin_RID),
    .m_axi_gmem_cin_RUSER(m_axi_gmem_cin_RUSER),
    .m_axi_gmem_cin_RRESP(m_axi_gmem_cin_RRESP),
    .m_axi_gmem_cin_BVALID(m_axi_gmem_cin_BVALID),
    .m_axi_gmem_cin_BREADY(m_axi_gmem_cin_BREADY),
    .m_axi_gmem_cin_BRESP(m_axi_gmem_cin_BRESP),
    .m_axi_gmem_cin_BID(m_axi_gmem_cin_BID),
    .m_axi_gmem_cin_BUSER(m_axi_gmem_cin_BUSER),
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start_Boundary_X4Y2_To_X6Y2(ap_start_Boundary_X4Y2_To_X6Y2_out),
    .ap_rst_n_Boundary_X4Y2_To_X6Y2(ap_rst_n_Boundary_X4Y2_To_X6Y2_out),
    .ap_done_Boundary_X4Y2_To_X6Y2(ap_done_Boundary_X4Y2_To_X6Y2_in),
    .ap_start_Boundary_X6Y0_To_X6Y2(ap_start_Boundary_X6Y0_To_X6Y2_out),
    .ap_rst_n_Boundary_X6Y0_To_X6Y2(ap_rst_n_Boundary_X6Y0_To_X6Y2_out),
    .ap_done_Boundary_X6Y0_To_X6Y2(ap_done_Boundary_X6Y0_To_X6Y2_in),
    .ap_start_Boundary_X4Y0_To_X4Y2(ap_start_Boundary_X4Y0_To_X4Y2_out),
    .ap_rst_n_Boundary_X4Y0_To_X4Y2(ap_rst_n_Boundary_X4Y0_To_X4Y2_out),
    .ap_done_Boundary_X4Y0_To_X4Y2(ap_done_Boundary_X4Y0_To_X4Y2_in)
  );


  (* keep_hierarchy = "yes" *) CR_X4Y4_To_CR_X5Y5_ctrl CR_X4Y4_To_CR_X5Y5_ctrl_U0 (
    .PE_wrapper190_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper190_U0_fifo_w_out_V_V_din_pass_0_in),
    .PE_wrapper190_U0_fifo_w_out_V_V_din_pass_1(PE_wrapper190_U0_fifo_w_out_V_V_din_pass_1_out),
    .fifo_w_PE_3_5_V_V_full_n_pass_0(fifo_w_PE_3_5_V_V_full_n_pass_0_out),
    .fifo_w_PE_3_5_V_V_full_n_pass_1(fifo_w_PE_3_5_V_V_full_n_pass_1_in),
    .PE_wrapper190_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper190_U0_fifo_w_out_V_V_write_pass_0_in),
    .PE_wrapper190_U0_fifo_w_out_V_V_write_pass_1(PE_wrapper190_U0_fifo_w_out_V_V_write_pass_1_out),
    .PE_wrapper179_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper179_U0_fifo_cin_out_V_V_din_pass_0_in),
    .PE_wrapper179_U0_fifo_cin_out_V_V_din_pass_1(PE_wrapper179_U0_fifo_cin_out_V_V_din_pass_1_out),
    .fifo_cin_PE_3_5_V_V_full_n_pass_0(fifo_cin_PE_3_5_V_V_full_n_pass_0_out),
    .fifo_cin_PE_3_5_V_V_full_n_pass_1(fifo_cin_PE_3_5_V_V_full_n_pass_1_in),
    .PE_wrapper179_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper179_U0_fifo_cin_out_V_V_write_pass_0_in),
    .PE_wrapper179_U0_fifo_cin_out_V_V_write_pass_1(PE_wrapper179_U0_fifo_cin_out_V_V_write_pass_1_out),
    .kernel0_entry12_U0_cout_V_out_din_pass_1(kernel0_entry12_U0_cout_V_out_din_pass_1_in),
    .kernel0_entry12_U0_cout_V_out_din_pass_2(kernel0_entry12_U0_cout_V_out_din_pass_2_out),
    .cout_V_c_full_n_pass_1(cout_V_c_full_n_pass_1_out),
    .cout_V_c_full_n_pass_2(cout_V_c_full_n_pass_2_in),
    .kernel0_entry12_U0_cout_V_out_write_pass_1(kernel0_entry12_U0_cout_V_out_write_pass_1_in),
    .kernel0_entry12_U0_cout_V_out_write_pass_2(kernel0_entry12_U0_cout_V_out_write_pass_2_out),
    .PE_wrapper190_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper190_U0_fifo_cin_out_V_V_din_pass_0_in),
    .fifo_cin_PE_4_4_V_V_full_n_pass_0(fifo_cin_PE_4_4_V_V_full_n_pass_0_out),
    .PE_wrapper190_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper190_U0_fifo_cin_out_V_V_write_pass_0_in),
    .PE_wrapper201_U0_fifo_w_out_V_V_din_pass_1(PE_wrapper201_U0_fifo_w_out_V_V_din_pass_1_in),
    .fifo_w_PE_4_4_V_V_full_n_pass_1(fifo_w_PE_4_4_V_V_full_n_pass_1_out),
    .PE_wrapper201_U0_fifo_w_out_V_V_write_pass_1(PE_wrapper201_U0_fifo_w_out_V_V_write_pass_1_in),
    .cout_drain_IO_L1_out_wrapper440_U0_fifo_cout_drain_out_V_V_din_pass_1(cout_drain_IO_L1_out_wrapper440_U0_fifo_cout_drain_out_V_V_din_pass_1_in),
    .fifo_cout_drain_cout_drain_IO_L1_out_4_6_V_V_full_n_pass_1(fifo_cout_drain_cout_drain_IO_L1_out_4_6_V_V_full_n_pass_1_out),
    .cout_drain_IO_L1_out_wrapper440_U0_fifo_cout_drain_out_V_V_write_pass_1(cout_drain_IO_L1_out_wrapper440_U0_fifo_cout_drain_out_V_V_write_pass_1_in),
    .PE_wrapper213_U0_fifo_w_out_V_V_din_pass_2(PE_wrapper213_U0_fifo_w_out_V_V_din_pass_2_in),
    .fifo_w_PE_5_4_V_V_full_n_pass_2(fifo_w_PE_5_4_V_V_full_n_pass_2_out),
    .PE_wrapper213_U0_fifo_w_out_V_V_write_pass_2(PE_wrapper213_U0_fifo_w_out_V_V_write_pass_2_in),
    .PE_wrapper214_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper214_U0_fifo_w_out_V_V_din_pass_0_out),
    .fifo_w_PE_5_5_V_V_full_n_pass_0(fifo_w_PE_5_5_V_V_full_n_pass_0_in),
    .PE_wrapper214_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper214_U0_fifo_w_out_V_V_write_pass_0_out),
    .cout_drain_IO_L1_out_wrapper441_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper441_U0_fifo_cout_drain_out_V_V_din_pass_0_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_4_5_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_4_5_V_V_full_n_pass_0_in),
    .cout_drain_IO_L1_out_wrapper441_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper441_U0_fifo_cout_drain_out_V_V_write_pass_0_out),
    .w_IO_L3_in_serialize_U0_fifo_w_local_out_V_V_din_pass_0(w_IO_L3_in_serialize_U0_fifo_w_local_out_V_V_din_pass_0_out),
    .fifo_w_w_IO_L3_in_serialize_V_V_full_n_pass_0(fifo_w_w_IO_L3_in_serialize_V_V_full_n_pass_0_in),
    .w_IO_L3_in_serialize_U0_fifo_w_local_out_V_V_write_pass_0(w_IO_L3_in_serialize_U0_fifo_w_local_out_V_V_write_pass_0_out),
    .PE_wrapper214_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper214_U0_fifo_cin_out_V_V_din_pass_0_out),
    .fifo_cin_PE_6_4_V_V_full_n_pass_0(fifo_cin_PE_6_4_V_V_full_n_pass_0_in),
    .PE_wrapper214_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper214_U0_fifo_cin_out_V_V_write_pass_0_out),
    .PE_wrapper202_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper202_U0_fifo_w_out_V_V_din_pass_0_out),
    .fifo_w_PE_4_5_V_V_full_n_pass_0(fifo_w_PE_4_5_V_V_full_n_pass_0_in),
    .PE_wrapper202_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper202_U0_fifo_w_out_V_V_write_pass_0_out),
    .PE_wrapper202_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper202_U0_fifo_cout_drain_out_V_din_pass_0_out),
    .fifo_cout_drain_PE_4_4_V_full_n_pass_0(fifo_cout_drain_PE_4_4_V_full_n_pass_0_in),
    .PE_wrapper202_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper202_U0_fifo_cout_drain_out_V_write_pass_0_out),
    .kernel0_entry12_U0_w_V_out_din_pass_1(kernel0_entry12_U0_w_V_out_din_pass_1_in),
    .w_V_c_full_n_pass_1(w_V_c_full_n_pass_1_out),
    .kernel0_entry12_U0_w_V_out_write_pass_1(kernel0_entry12_U0_w_V_out_write_pass_1_in),
    .m_axi_gmem_w_AWVALID(m_axi_gmem_w_AWVALID),
    .m_axi_gmem_w_AWREADY(m_axi_gmem_w_AWREADY),
    .m_axi_gmem_w_AWADDR(m_axi_gmem_w_AWADDR),
    .m_axi_gmem_w_AWID(m_axi_gmem_w_AWID),
    .m_axi_gmem_w_AWLEN(m_axi_gmem_w_AWLEN),
    .m_axi_gmem_w_AWSIZE(m_axi_gmem_w_AWSIZE),
    .m_axi_gmem_w_AWBURST(m_axi_gmem_w_AWBURST),
    .m_axi_gmem_w_AWLOCK(m_axi_gmem_w_AWLOCK),
    .m_axi_gmem_w_AWCACHE(m_axi_gmem_w_AWCACHE),
    .m_axi_gmem_w_AWPROT(m_axi_gmem_w_AWPROT),
    .m_axi_gmem_w_AWQOS(m_axi_gmem_w_AWQOS),
    .m_axi_gmem_w_AWREGION(m_axi_gmem_w_AWREGION),
    .m_axi_gmem_w_AWUSER(m_axi_gmem_w_AWUSER),
    .m_axi_gmem_w_WVALID(m_axi_gmem_w_WVALID),
    .m_axi_gmem_w_WREADY(m_axi_gmem_w_WREADY),
    .m_axi_gmem_w_WDATA(m_axi_gmem_w_WDATA),
    .m_axi_gmem_w_WSTRB(m_axi_gmem_w_WSTRB),
    .m_axi_gmem_w_WLAST(m_axi_gmem_w_WLAST),
    .m_axi_gmem_w_WID(m_axi_gmem_w_WID),
    .m_axi_gmem_w_WUSER(m_axi_gmem_w_WUSER),
    .m_axi_gmem_w_ARVALID(m_axi_gmem_w_ARVALID),
    .m_axi_gmem_w_ARREADY(m_axi_gmem_w_ARREADY),
    .m_axi_gmem_w_ARADDR(m_axi_gmem_w_ARADDR),
    .m_axi_gmem_w_ARID(m_axi_gmem_w_ARID),
    .m_axi_gmem_w_ARLEN(m_axi_gmem_w_ARLEN),
    .m_axi_gmem_w_ARSIZE(m_axi_gmem_w_ARSIZE),
    .m_axi_gmem_w_ARBURST(m_axi_gmem_w_ARBURST),
    .m_axi_gmem_w_ARLOCK(m_axi_gmem_w_ARLOCK),
    .m_axi_gmem_w_ARCACHE(m_axi_gmem_w_ARCACHE),
    .m_axi_gmem_w_ARPROT(m_axi_gmem_w_ARPROT),
    .m_axi_gmem_w_ARQOS(m_axi_gmem_w_ARQOS),
    .m_axi_gmem_w_ARREGION(m_axi_gmem_w_ARREGION),
    .m_axi_gmem_w_ARUSER(m_axi_gmem_w_ARUSER),
    .m_axi_gmem_w_RVALID(m_axi_gmem_w_RVALID),
    .m_axi_gmem_w_RREADY(m_axi_gmem_w_RREADY),
    .m_axi_gmem_w_RDATA(m_axi_gmem_w_RDATA),
    .m_axi_gmem_w_RLAST(m_axi_gmem_w_RLAST),
    .m_axi_gmem_w_RID(m_axi_gmem_w_RID),
    .m_axi_gmem_w_RUSER(m_axi_gmem_w_RUSER),
    .m_axi_gmem_w_RRESP(m_axi_gmem_w_RRESP),
    .m_axi_gmem_w_BVALID(m_axi_gmem_w_BVALID),
    .m_axi_gmem_w_BREADY(m_axi_gmem_w_BREADY),
    .m_axi_gmem_w_BRESP(m_axi_gmem_w_BRESP),
    .m_axi_gmem_w_BID(m_axi_gmem_w_BID),
    .m_axi_gmem_w_BUSER(m_axi_gmem_w_BUSER),
    .ap_clk(ap_clk),
    .ap_start_Boundary_X4Y4_To_X6Y4(ap_start_Boundary_X4Y4_To_X6Y4_in),
    .ap_rst_n_Boundary_X4Y4_To_X6Y4(ap_rst_n_Boundary_X4Y4_To_X6Y4_in),
    .ap_done_Boundary_X4Y4_To_X6Y4(ap_done_Boundary_X4Y4_To_X6Y4_out),
    .ap_start_Boundary_X4Y6_To_X6Y6(ap_start_Boundary_X4Y6_To_X6Y6_out),
    .ap_rst_n_Boundary_X4Y6_To_X6Y6(ap_rst_n_Boundary_X4Y6_To_X6Y6_out),
    .ap_done_Boundary_X4Y6_To_X6Y6(ap_done_Boundary_X4Y6_To_X6Y6_in)
  );


  (* keep_hierarchy = "yes" *) CR_X4Y12_To_CR_X5Y13_ctrl CR_X4Y12_To_CR_X5Y13_ctrl_U0 (
    .PE_wrapper230_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper230_U0_fifo_w_out_V_V_din_pass_0_in),
    .PE_wrapper230_U0_fifo_w_out_V_V_din_pass_1(PE_wrapper230_U0_fifo_w_out_V_V_din_pass_1_out),
    .fifo_w_PE_6_9_V_V_full_n_pass_0(fifo_w_PE_6_9_V_V_full_n_pass_0_out),
    .fifo_w_PE_6_9_V_V_full_n_pass_1(fifo_w_PE_6_9_V_V_full_n_pass_1_in),
    .PE_wrapper230_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper230_U0_fifo_w_out_V_V_write_pass_0_in),
    .PE_wrapper230_U0_fifo_w_out_V_V_write_pass_1(PE_wrapper230_U0_fifo_w_out_V_V_write_pass_1_out),
    .cout_drain_IO_L1_out_wrapper522_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper522_U0_fifo_cout_drain_out_V_V_din_pass_0_in),
    .cout_drain_IO_L1_out_wrapper522_U0_fifo_cout_drain_out_V_V_din_pass_1(cout_drain_IO_L1_out_wrapper522_U0_fifo_cout_drain_out_V_V_din_pass_1_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_9_4_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_9_4_V_V_full_n_pass_0_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_9_4_V_V_full_n_pass_1(fifo_cout_drain_cout_drain_IO_L1_out_9_4_V_V_full_n_pass_1_in),
    .cout_drain_IO_L1_out_wrapper522_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper522_U0_fifo_cout_drain_out_V_V_write_pass_0_in),
    .cout_drain_IO_L1_out_wrapper522_U0_fifo_cout_drain_out_V_V_write_pass_1(cout_drain_IO_L1_out_wrapper522_U0_fifo_cout_drain_out_V_V_write_pass_1_out),
    .cout_drain_IO_L1_out_wrapper542_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper542_U0_fifo_cout_drain_out_V_V_din_pass_0_in),
    .cout_drain_IO_L1_out_wrapper542_U0_fifo_cout_drain_out_V_V_din_pass_1(cout_drain_IO_L1_out_wrapper542_U0_fifo_cout_drain_out_V_V_din_pass_1_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_10_0_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_10_0_V_V_full_n_pass_0_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_10_0_V_V_full_n_pass_1(fifo_cout_drain_cout_drain_IO_L1_out_10_0_V_V_full_n_pass_1_in),
    .cout_drain_IO_L1_out_wrapper542_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper542_U0_fifo_cout_drain_out_V_V_write_pass_0_in),
    .cout_drain_IO_L1_out_wrapper542_U0_fifo_cout_drain_out_V_V_write_pass_1(cout_drain_IO_L1_out_wrapper542_U0_fifo_cout_drain_out_V_V_write_pass_1_out),
    .PE_wrapper219_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper219_U0_fifo_cin_out_V_V_din_pass_0_in),
    .PE_wrapper219_U0_fifo_cin_out_V_V_din_pass_1(PE_wrapper219_U0_fifo_cin_out_V_V_din_pass_1_out),
    .fifo_cin_PE_6_9_V_V_full_n_pass_0(fifo_cin_PE_6_9_V_V_full_n_pass_0_out),
    .fifo_cin_PE_6_9_V_V_full_n_pass_1(fifo_cin_PE_6_9_V_V_full_n_pass_1_in),
    .PE_wrapper219_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper219_U0_fifo_cin_out_V_V_write_pass_0_in),
    .PE_wrapper219_U0_fifo_cin_out_V_V_write_pass_1(PE_wrapper219_U0_fifo_cin_out_V_V_write_pass_1_out),
    .PE_wrapper172_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper172_U0_fifo_cin_out_V_V_din_pass_0_in),
    .PE_wrapper172_U0_fifo_cin_out_V_V_din_pass_1(PE_wrapper172_U0_fifo_cin_out_V_V_din_pass_1_out),
    .fifo_cin_PE_2_10_V_V_full_n_pass_0(fifo_cin_PE_2_10_V_V_full_n_pass_0_out),
    .fifo_cin_PE_2_10_V_V_full_n_pass_1(fifo_cin_PE_2_10_V_V_full_n_pass_1_in),
    .PE_wrapper172_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper172_U0_fifo_cin_out_V_V_write_pass_0_in),
    .PE_wrapper172_U0_fifo_cin_out_V_V_write_pass_1(PE_wrapper172_U0_fifo_cin_out_V_V_write_pass_1_out),
    .cin_IO_L2_in134_U0_fifo_cin_out_V_V_din_pass_0(cin_IO_L2_in134_U0_fifo_cin_out_V_V_din_pass_0_in),
    .cin_IO_L2_in134_U0_fifo_cin_out_V_V_din_pass_1(cin_IO_L2_in134_U0_fifo_cin_out_V_V_din_pass_1_out),
    .fifo_cin_cin_IO_L2_in_11_V_V_full_n_pass_0(fifo_cin_cin_IO_L2_in_11_V_V_full_n_pass_0_out),
    .fifo_cin_cin_IO_L2_in_11_V_V_full_n_pass_1(fifo_cin_cin_IO_L2_in_11_V_V_full_n_pass_1_in),
    .cin_IO_L2_in134_U0_fifo_cin_out_V_V_write_pass_0(cin_IO_L2_in134_U0_fifo_cin_out_V_V_write_pass_0_in),
    .cin_IO_L2_in134_U0_fifo_cin_out_V_V_write_pass_1(cin_IO_L2_in134_U0_fifo_cin_out_V_V_write_pass_1_out),
    .PE_wrapper194_U0_fifo_w_out_V_V_din_pass_1(PE_wrapper194_U0_fifo_w_out_V_V_din_pass_1_in),
    .PE_wrapper194_U0_fifo_w_out_V_V_din_pass_2(PE_wrapper194_U0_fifo_w_out_V_V_din_pass_2_out),
    .fifo_w_PE_3_9_V_V_full_n_pass_1(fifo_w_PE_3_9_V_V_full_n_pass_1_out),
    .fifo_w_PE_3_9_V_V_full_n_pass_2(fifo_w_PE_3_9_V_V_full_n_pass_2_in),
    .PE_wrapper194_U0_fifo_w_out_V_V_write_pass_1(PE_wrapper194_U0_fifo_w_out_V_V_write_pass_1_in),
    .PE_wrapper194_U0_fifo_w_out_V_V_write_pass_2(PE_wrapper194_U0_fifo_w_out_V_V_write_pass_2_out),
    .cout_drain_IO_L1_out_wrapper548_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper548_U0_fifo_cout_drain_out_V_V_din_pass_0_in),
    .cout_drain_IO_L1_out_wrapper548_U0_fifo_cout_drain_out_V_V_din_pass_1(cout_drain_IO_L1_out_wrapper548_U0_fifo_cout_drain_out_V_V_din_pass_1_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_11_9_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_11_9_V_V_full_n_pass_0_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_11_9_V_V_full_n_pass_1(fifo_cout_drain_cout_drain_IO_L1_out_11_9_V_V_full_n_pass_1_in),
    .cout_drain_IO_L1_out_wrapper548_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper548_U0_fifo_cout_drain_out_V_V_write_pass_0_in),
    .cout_drain_IO_L1_out_wrapper548_U0_fifo_cout_drain_out_V_V_write_pass_1(cout_drain_IO_L1_out_wrapper548_U0_fifo_cout_drain_out_V_V_write_pass_1_out),
    .PE_wrapper219_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper219_U0_fifo_cout_drain_out_V_din_pass_0_in),
    .PE_wrapper219_U0_fifo_cout_drain_out_V_din_pass_1(PE_wrapper219_U0_fifo_cout_drain_out_V_din_pass_1_out),
    .fifo_cout_drain_PE_5_9_V_full_n_pass_0(fifo_cout_drain_PE_5_9_V_full_n_pass_0_out),
    .fifo_cout_drain_PE_5_9_V_full_n_pass_1(fifo_cout_drain_PE_5_9_V_full_n_pass_1_in),
    .PE_wrapper219_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper219_U0_fifo_cout_drain_out_V_write_pass_0_in),
    .PE_wrapper219_U0_fifo_cout_drain_out_V_write_pass_1(PE_wrapper219_U0_fifo_cout_drain_out_V_write_pass_1_out),
    .cout_drain_IO_L1_out_wrapper517_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper517_U0_fifo_cout_drain_out_V_V_din_pass_0_in),
    .cout_drain_IO_L1_out_wrapper517_U0_fifo_cout_drain_out_V_V_din_pass_1(cout_drain_IO_L1_out_wrapper517_U0_fifo_cout_drain_out_V_V_din_pass_1_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_9_9_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_9_9_V_V_full_n_pass_0_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_9_9_V_V_full_n_pass_1(fifo_cout_drain_cout_drain_IO_L1_out_9_9_V_V_full_n_pass_1_in),
    .cout_drain_IO_L1_out_wrapper517_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper517_U0_fifo_cout_drain_out_V_V_write_pass_0_in),
    .cout_drain_IO_L1_out_wrapper517_U0_fifo_cout_drain_out_V_V_write_pass_1(cout_drain_IO_L1_out_wrapper517_U0_fifo_cout_drain_out_V_V_write_pass_1_out),
    .cout_drain_IO_L1_out_wrapper533_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper533_U0_fifo_cout_drain_out_V_V_din_pass_0_in),
    .cout_drain_IO_L1_out_wrapper533_U0_fifo_cout_drain_out_V_V_din_pass_1(cout_drain_IO_L1_out_wrapper533_U0_fifo_cout_drain_out_V_V_din_pass_1_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_10_9_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_10_9_V_V_full_n_pass_0_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_10_9_V_V_full_n_pass_1(fifo_cout_drain_cout_drain_IO_L1_out_10_9_V_V_full_n_pass_1_in),
    .cout_drain_IO_L1_out_wrapper533_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper533_U0_fifo_cout_drain_out_V_V_write_pass_0_in),
    .cout_drain_IO_L1_out_wrapper533_U0_fifo_cout_drain_out_V_V_write_pass_1(cout_drain_IO_L1_out_wrapper533_U0_fifo_cout_drain_out_V_V_write_pass_1_out),
    .cout_drain_IO_L1_out_wrapper535_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper535_U0_fifo_cout_drain_out_V_V_din_pass_0_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_10_7_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_10_7_V_V_full_n_pass_0_in),
    .cout_drain_IO_L1_out_wrapper535_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper535_U0_fifo_cout_drain_out_V_V_write_pass_0_out),
    .PE_wrapper219_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper219_U0_fifo_w_out_V_V_din_pass_0_in),
    .fifo_w_PE_5_10_V_V_full_n_pass_0(fifo_w_PE_5_10_V_V_full_n_pass_0_out),
    .PE_wrapper219_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper219_U0_fifo_w_out_V_V_write_pass_0_in),
    .cout_drain_IO_L1_out_wrapper537_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper537_U0_fifo_cout_drain_out_V_V_din_pass_0_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_10_5_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_10_5_V_V_full_n_pass_0_in),
    .cout_drain_IO_L1_out_wrapper537_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper537_U0_fifo_cout_drain_out_V_V_write_pass_0_out),
    .PE_wrapper171_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper171_U0_fifo_cin_out_V_V_din_pass_0_in),
    .fifo_cin_PE_2_9_V_V_full_n_pass_0(fifo_cin_PE_2_9_V_V_full_n_pass_0_out),
    .PE_wrapper171_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper171_U0_fifo_cin_out_V_V_write_pass_0_in),
    .PE_wrapper172_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper172_U0_fifo_w_out_V_V_din_pass_0_in),
    .fifo_w_PE_1_11_V_V_full_n_pass_0(fifo_w_PE_1_11_V_V_full_n_pass_0_out),
    .PE_wrapper172_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper172_U0_fifo_w_out_V_V_write_pass_0_in),
    .cout_drain_IO_L1_out_wrapper551_U0_fifo_cout_drain_out_V_V_din_pass_1(cout_drain_IO_L1_out_wrapper551_U0_fifo_cout_drain_out_V_V_din_pass_1_in),
    .fifo_cout_drain_cout_drain_IO_L1_out_11_6_V_V_full_n_pass_1(fifo_cout_drain_cout_drain_IO_L1_out_11_6_V_V_full_n_pass_1_out),
    .cout_drain_IO_L1_out_wrapper551_U0_fifo_cout_drain_out_V_V_write_pass_1(cout_drain_IO_L1_out_wrapper551_U0_fifo_cout_drain_out_V_V_write_pass_1_in),
    .cout_drain_IO_L1_out_wrapper555_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper555_U0_fifo_cout_drain_out_V_V_din_pass_0_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_11_2_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_11_2_V_V_full_n_pass_0_in),
    .cout_drain_IO_L1_out_wrapper555_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper555_U0_fifo_cout_drain_out_V_V_write_pass_0_out),
    .PE_wrapper196_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper196_U0_fifo_cin_out_V_V_din_pass_0_in),
    .fifo_cin_PE_4_10_V_V_full_n_pass_0(fifo_cin_PE_4_10_V_V_full_n_pass_0_out),
    .PE_wrapper196_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper196_U0_fifo_cin_out_V_V_write_pass_0_in),
    .cout_drain_IO_L1_out_wrapper539_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper539_U0_fifo_cout_drain_out_V_V_din_pass_0_in),
    .fifo_cout_drain_cout_drain_IO_L1_out_10_3_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_10_3_V_V_full_n_pass_0_out),
    .cout_drain_IO_L1_out_wrapper539_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper539_U0_fifo_cout_drain_out_V_V_write_pass_0_in),
    .PE_wrapper244_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper244_U0_fifo_cin_out_V_V_din_pass_0_out),
    .fifo_cin_PE_8_10_V_V_full_n_pass_0(fifo_cin_PE_8_10_V_V_full_n_pass_0_in),
    .PE_wrapper244_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper244_U0_fifo_cin_out_V_V_write_pass_0_out),
    .PE_wrapper231_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper231_U0_fifo_w_out_V_V_din_pass_0_in),
    .fifo_w_PE_6_10_V_V_full_n_pass_0(fifo_w_PE_6_10_V_V_full_n_pass_0_out),
    .PE_wrapper231_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper231_U0_fifo_w_out_V_V_write_pass_0_in),
    .PE_wrapper173_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper173_U0_fifo_w_out_V_V_din_pass_0_out),
    .fifo_w_PE_1_12_V_V_full_n_pass_0(fifo_w_PE_1_12_V_V_full_n_pass_0_in),
    .PE_wrapper173_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper173_U0_fifo_w_out_V_V_write_pass_0_out),
    .PE_wrapper231_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper231_U0_fifo_cout_drain_out_V_din_pass_0_in),
    .fifo_cout_drain_PE_6_9_V_full_n_pass_0(fifo_cout_drain_PE_6_9_V_full_n_pass_0_out),
    .PE_wrapper231_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper231_U0_fifo_cout_drain_out_V_write_pass_0_in),
    .PE_wrapper207_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper207_U0_fifo_w_out_V_V_din_pass_0_in),
    .fifo_w_PE_4_10_V_V_full_n_pass_0(fifo_w_PE_4_10_V_V_full_n_pass_0_out),
    .PE_wrapper207_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper207_U0_fifo_w_out_V_V_write_pass_0_in),
    .PE_wrapper221_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper221_U0_fifo_cout_drain_out_V_din_pass_0_in),
    .fifo_cout_drain_PE_5_11_V_full_n_pass_0(fifo_cout_drain_PE_5_11_V_full_n_pass_0_out),
    .PE_wrapper221_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper221_U0_fifo_cout_drain_out_V_write_pass_0_in),
    .PE_wrapper183_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper183_U0_fifo_cout_drain_out_V_din_pass_0_out),
    .fifo_cout_drain_PE_2_9_V_full_n_pass_0(fifo_cout_drain_PE_2_9_V_full_n_pass_0_in),
    .PE_wrapper183_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper183_U0_fifo_cout_drain_out_V_write_pass_0_out),
    .PE_wrapper161_U0_fifo_cin_out_V_V_din_pass_1(PE_wrapper161_U0_fifo_cin_out_V_V_din_pass_1_in),
    .fifo_cin_PE_1_11_V_V_full_n_pass_1(fifo_cin_PE_1_11_V_V_full_n_pass_1_out),
    .PE_wrapper161_U0_fifo_cin_out_V_V_write_pass_1(PE_wrapper161_U0_fifo_cin_out_V_V_write_pass_1_in),
    .PE_wrapper232_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper232_U0_fifo_cout_drain_out_V_din_pass_0_out),
    .fifo_cout_drain_PE_6_10_V_full_n_pass_0(fifo_cout_drain_PE_6_10_V_full_n_pass_0_in),
    .PE_wrapper232_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper232_U0_fifo_cout_drain_out_V_write_pass_0_out),
    .kernel0_entry12_U0_cout_V_out_din_pass_5(kernel0_entry12_U0_cout_V_out_din_pass_5_in),
    .cout_V_c_full_n_pass_5(cout_V_c_full_n_pass_5_out),
    .kernel0_entry12_U0_cout_V_out_write_pass_5(kernel0_entry12_U0_cout_V_out_write_pass_5_in),
    .cout_drain_IO_L1_out_wrapper540_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper540_U0_fifo_cout_drain_out_V_V_din_pass_0_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_10_2_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_10_2_V_V_full_n_pass_0_in),
    .cout_drain_IO_L1_out_wrapper540_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper540_U0_fifo_cout_drain_out_V_V_write_pass_0_out),
    .cout_drain_IO_L1_out_wrapper552_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper552_U0_fifo_cout_drain_out_V_V_din_pass_0_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_11_5_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_11_5_V_V_full_n_pass_0_in),
    .cout_drain_IO_L1_out_wrapper552_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper552_U0_fifo_cout_drain_out_V_V_write_pass_0_out),
    .PE_wrapper243_U0_fifo_w_out_V_V_din_pass_3(PE_wrapper243_U0_fifo_w_out_V_V_din_pass_3_in),
    .fifo_w_PE_7_10_V_V_full_n_pass_3(fifo_w_PE_7_10_V_V_full_n_pass_3_out),
    .PE_wrapper243_U0_fifo_w_out_V_V_write_pass_3(PE_wrapper243_U0_fifo_w_out_V_V_write_pass_3_in),
    .PE_wrapper243_U0_fifo_cout_drain_out_V_din_pass_3(PE_wrapper243_U0_fifo_cout_drain_out_V_din_pass_3_in),
    .fifo_cout_drain_PE_7_9_V_full_n_pass_3(fifo_cout_drain_PE_7_9_V_full_n_pass_3_out),
    .PE_wrapper243_U0_fifo_cout_drain_out_V_write_pass_3(PE_wrapper243_U0_fifo_cout_drain_out_V_write_pass_3_in),
    .PE_wrapper184_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper184_U0_fifo_cout_drain_out_V_din_pass_0_in),
    .fifo_cout_drain_PE_2_10_V_full_n_pass_0(fifo_cout_drain_PE_2_10_V_full_n_pass_0_out),
    .PE_wrapper184_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper184_U0_fifo_cout_drain_out_V_write_pass_0_in),
    .PE_wrapper243_U0_fifo_cin_out_V_V_din_pass_3(PE_wrapper243_U0_fifo_cin_out_V_V_din_pass_3_in),
    .fifo_cin_PE_8_9_V_V_full_n_pass_3(fifo_cin_PE_8_9_V_V_full_n_pass_3_out),
    .PE_wrapper243_U0_fifo_cin_out_V_V_write_pass_3(PE_wrapper243_U0_fifo_cin_out_V_V_write_pass_3_in),
    .PE_wrapper255_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper255_U0_fifo_cout_drain_out_V_din_pass_0_out),
    .fifo_cout_drain_PE_8_9_V_full_n_pass_0(fifo_cout_drain_PE_8_9_V_full_n_pass_0_in),
    .PE_wrapper255_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper255_U0_fifo_cout_drain_out_V_write_pass_0_out),
    .PE_wrapper185_U0_fifo_cout_drain_out_V_din_pass_1(PE_wrapper185_U0_fifo_cout_drain_out_V_din_pass_1_in),
    .fifo_cout_drain_PE_2_11_V_full_n_pass_1(fifo_cout_drain_PE_2_11_V_full_n_pass_1_out),
    .PE_wrapper185_U0_fifo_cout_drain_out_V_write_pass_1(PE_wrapper185_U0_fifo_cout_drain_out_V_write_pass_1_in),
    .cout_drain_IO_L1_out_wrapper518_U0_fifo_cout_drain_out_V_V_din_pass_1(cout_drain_IO_L1_out_wrapper518_U0_fifo_cout_drain_out_V_V_din_pass_1_in),
    .fifo_cout_drain_cout_drain_IO_L1_out_9_8_V_V_full_n_pass_1(fifo_cout_drain_cout_drain_IO_L1_out_9_8_V_V_full_n_pass_1_out),
    .cout_drain_IO_L1_out_wrapper518_U0_fifo_cout_drain_out_V_V_write_pass_1(cout_drain_IO_L1_out_wrapper518_U0_fifo_cout_drain_out_V_V_write_pass_1_in),
    .PE_wrapper255_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper255_U0_fifo_cin_out_V_V_din_pass_0_out),
    .fifo_cin_PE_9_9_V_V_full_n_pass_0(fifo_cin_PE_9_9_V_V_full_n_pass_0_in),
    .PE_wrapper255_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper255_U0_fifo_cin_out_V_V_write_pass_0_out),
    .PE_wrapper244_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper244_U0_fifo_w_out_V_V_din_pass_0_out),
    .fifo_w_PE_7_11_V_V_full_n_pass_0(fifo_w_PE_7_11_V_V_full_n_pass_0_in),
    .PE_wrapper244_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper244_U0_fifo_w_out_V_V_write_pass_0_out),
    .PE_wrapper173_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper173_U0_fifo_cout_drain_out_V_din_pass_0_out),
    .fifo_cout_drain_PE_1_11_V_full_n_pass_0(fifo_cout_drain_PE_1_11_V_full_n_pass_0_in),
    .PE_wrapper173_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper173_U0_fifo_cout_drain_out_V_write_pass_0_out),
    .PE_wrapper254_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper254_U0_fifo_w_out_V_V_din_pass_0_in),
    .fifo_w_PE_8_9_V_V_full_n_pass_0(fifo_w_PE_8_9_V_V_full_n_pass_0_out),
    .PE_wrapper254_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper254_U0_fifo_w_out_V_V_write_pass_0_in),
    .PE_wrapper208_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper208_U0_fifo_cout_drain_out_V_din_pass_0_out),
    .fifo_cout_drain_PE_4_10_V_full_n_pass_0(fifo_cout_drain_PE_4_10_V_full_n_pass_0_in),
    .PE_wrapper208_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper208_U0_fifo_cout_drain_out_V_write_pass_0_out),
    .cout_drain_IO_L1_out_wrapper536_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper536_U0_fifo_cout_drain_out_V_V_din_pass_0_in),
    .fifo_cout_drain_cout_drain_IO_L1_out_10_6_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_10_6_V_V_full_n_pass_0_out),
    .cout_drain_IO_L1_out_wrapper536_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper536_U0_fifo_cout_drain_out_V_V_write_pass_0_in),
    .PE_wrapper182_U0_fifo_w_out_V_V_din_pass_1(PE_wrapper182_U0_fifo_w_out_V_V_din_pass_1_in),
    .fifo_w_PE_2_9_V_V_full_n_pass_1(fifo_w_PE_2_9_V_V_full_n_pass_1_out),
    .PE_wrapper182_U0_fifo_w_out_V_V_write_pass_1(PE_wrapper182_U0_fifo_w_out_V_V_write_pass_1_in),
    .PE_wrapper220_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper220_U0_fifo_w_out_V_V_din_pass_0_out),
    .fifo_w_PE_5_11_V_V_full_n_pass_0(fifo_w_PE_5_11_V_V_full_n_pass_0_in),
    .PE_wrapper220_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper220_U0_fifo_w_out_V_V_write_pass_0_out),
    .PE_wrapper255_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper255_U0_fifo_w_out_V_V_din_pass_0_out),
    .fifo_w_PE_8_10_V_V_full_n_pass_0(fifo_w_PE_8_10_V_V_full_n_pass_0_in),
    .PE_wrapper255_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper255_U0_fifo_w_out_V_V_write_pass_0_out),
    .cout_drain_IO_L1_out_wrapper534_U0_fifo_cout_drain_out_V_V_din_pass_1(cout_drain_IO_L1_out_wrapper534_U0_fifo_cout_drain_out_V_V_din_pass_1_in),
    .fifo_cout_drain_cout_drain_IO_L1_out_10_8_V_V_full_n_pass_1(fifo_cout_drain_cout_drain_IO_L1_out_10_8_V_V_full_n_pass_1_out),
    .cout_drain_IO_L1_out_wrapper534_U0_fifo_cout_drain_out_V_V_write_pass_1(cout_drain_IO_L1_out_wrapper534_U0_fifo_cout_drain_out_V_V_write_pass_1_in),
    .cout_drain_IO_L1_out_wrapper520_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper520_U0_fifo_cout_drain_out_V_V_din_pass_0_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_9_6_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_9_6_V_V_full_n_pass_0_in),
    .cout_drain_IO_L1_out_wrapper520_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper520_U0_fifo_cout_drain_out_V_V_write_pass_0_out),
    .cout_drain_IO_L3_out_U0_fifo_cout_drain_out_V_V_din_pass_2(cout_drain_IO_L3_out_U0_fifo_cout_drain_out_V_V_din_pass_2_in),
    .fifo_cout_drain_cout_drain_IO_L3_out_serialize_V_V_full_n_pass_2(fifo_cout_drain_cout_drain_IO_L3_out_serialize_V_V_full_n_pass_2_out),
    .cout_drain_IO_L3_out_U0_fifo_cout_drain_out_V_V_write_pass_2(cout_drain_IO_L3_out_U0_fifo_cout_drain_out_V_V_write_pass_2_in),
    .PE_wrapper173_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper173_U0_fifo_cin_out_V_V_din_pass_0_out),
    .fifo_cin_PE_2_11_V_V_full_n_pass_0(fifo_cin_PE_2_11_V_V_full_n_pass_0_in),
    .PE_wrapper173_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper173_U0_fifo_cin_out_V_V_write_pass_0_out),
    .PE_wrapper232_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper232_U0_fifo_w_out_V_V_din_pass_0_out),
    .fifo_w_PE_6_11_V_V_full_n_pass_0(fifo_w_PE_6_11_V_V_full_n_pass_0_in),
    .PE_wrapper232_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper232_U0_fifo_w_out_V_V_write_pass_0_out),
    .PE_wrapper183_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper183_U0_fifo_w_out_V_V_din_pass_0_out),
    .fifo_w_PE_2_10_V_V_full_n_pass_0(fifo_w_PE_2_10_V_V_full_n_pass_0_in),
    .PE_wrapper183_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper183_U0_fifo_w_out_V_V_write_pass_0_out),
    .PE_wrapper221_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper221_U0_fifo_w_out_V_V_din_pass_0_in),
    .fifo_w_PE_5_12_V_V_full_n_pass_0(fifo_w_PE_5_12_V_V_full_n_pass_0_out),
    .PE_wrapper221_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper221_U0_fifo_w_out_V_V_write_pass_0_in),
    .PE_wrapper208_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper208_U0_fifo_w_out_V_V_din_pass_0_out),
    .fifo_w_PE_4_11_V_V_full_n_pass_0(fifo_w_PE_4_11_V_V_full_n_pass_0_in),
    .PE_wrapper208_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper208_U0_fifo_w_out_V_V_write_pass_0_out),
    .PE_wrapper197_U0_fifo_cout_drain_out_V_din_pass_1(PE_wrapper197_U0_fifo_cout_drain_out_V_din_pass_1_in),
    .fifo_cout_drain_PE_3_11_V_full_n_pass_1(fifo_cout_drain_PE_3_11_V_full_n_pass_1_out),
    .PE_wrapper197_U0_fifo_cout_drain_out_V_write_pass_1(PE_wrapper197_U0_fifo_cout_drain_out_V_write_pass_1_in),
    .PE_wrapper183_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper183_U0_fifo_cin_out_V_V_din_pass_0_out),
    .fifo_cin_PE_3_9_V_V_full_n_pass_0(fifo_cin_PE_3_9_V_V_full_n_pass_0_in),
    .PE_wrapper183_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper183_U0_fifo_cin_out_V_V_write_pass_0_out),
    .cout_drain_IO_L1_out_wrapper553_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper553_U0_fifo_cout_drain_out_V_V_din_pass_0_in),
    .fifo_cout_drain_cout_drain_IO_L1_out_11_4_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_11_4_V_V_full_n_pass_0_out),
    .cout_drain_IO_L1_out_wrapper553_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper553_U0_fifo_cout_drain_out_V_V_write_pass_0_in),
    .m_axi_gmem_cout_AWVALID(m_axi_gmem_cout_AWVALID),
    .m_axi_gmem_cout_AWREADY(m_axi_gmem_cout_AWREADY),
    .m_axi_gmem_cout_AWADDR(m_axi_gmem_cout_AWADDR),
    .m_axi_gmem_cout_AWID(m_axi_gmem_cout_AWID),
    .m_axi_gmem_cout_AWLEN(m_axi_gmem_cout_AWLEN),
    .m_axi_gmem_cout_AWSIZE(m_axi_gmem_cout_AWSIZE),
    .m_axi_gmem_cout_AWBURST(m_axi_gmem_cout_AWBURST),
    .m_axi_gmem_cout_AWLOCK(m_axi_gmem_cout_AWLOCK),
    .m_axi_gmem_cout_AWCACHE(m_axi_gmem_cout_AWCACHE),
    .m_axi_gmem_cout_AWPROT(m_axi_gmem_cout_AWPROT),
    .m_axi_gmem_cout_AWQOS(m_axi_gmem_cout_AWQOS),
    .m_axi_gmem_cout_AWREGION(m_axi_gmem_cout_AWREGION),
    .m_axi_gmem_cout_AWUSER(m_axi_gmem_cout_AWUSER),
    .m_axi_gmem_cout_WVALID(m_axi_gmem_cout_WVALID),
    .m_axi_gmem_cout_WREADY(m_axi_gmem_cout_WREADY),
    .m_axi_gmem_cout_WDATA(m_axi_gmem_cout_WDATA),
    .m_axi_gmem_cout_WSTRB(m_axi_gmem_cout_WSTRB),
    .m_axi_gmem_cout_WLAST(m_axi_gmem_cout_WLAST),
    .m_axi_gmem_cout_WID(m_axi_gmem_cout_WID),
    .m_axi_gmem_cout_WUSER(m_axi_gmem_cout_WUSER),
    .m_axi_gmem_cout_ARVALID(m_axi_gmem_cout_ARVALID),
    .m_axi_gmem_cout_ARREADY(m_axi_gmem_cout_ARREADY),
    .m_axi_gmem_cout_ARADDR(m_axi_gmem_cout_ARADDR),
    .m_axi_gmem_cout_ARID(m_axi_gmem_cout_ARID),
    .m_axi_gmem_cout_ARLEN(m_axi_gmem_cout_ARLEN),
    .m_axi_gmem_cout_ARSIZE(m_axi_gmem_cout_ARSIZE),
    .m_axi_gmem_cout_ARBURST(m_axi_gmem_cout_ARBURST),
    .m_axi_gmem_cout_ARLOCK(m_axi_gmem_cout_ARLOCK),
    .m_axi_gmem_cout_ARCACHE(m_axi_gmem_cout_ARCACHE),
    .m_axi_gmem_cout_ARPROT(m_axi_gmem_cout_ARPROT),
    .m_axi_gmem_cout_ARQOS(m_axi_gmem_cout_ARQOS),
    .m_axi_gmem_cout_ARREGION(m_axi_gmem_cout_ARREGION),
    .m_axi_gmem_cout_ARUSER(m_axi_gmem_cout_ARUSER),
    .m_axi_gmem_cout_RVALID(m_axi_gmem_cout_RVALID),
    .m_axi_gmem_cout_RREADY(m_axi_gmem_cout_RREADY),
    .m_axi_gmem_cout_RDATA(m_axi_gmem_cout_RDATA),
    .m_axi_gmem_cout_RLAST(m_axi_gmem_cout_RLAST),
    .m_axi_gmem_cout_RID(m_axi_gmem_cout_RID),
    .m_axi_gmem_cout_RUSER(m_axi_gmem_cout_RUSER),
    .m_axi_gmem_cout_RRESP(m_axi_gmem_cout_RRESP),
    .m_axi_gmem_cout_BVALID(m_axi_gmem_cout_BVALID),
    .m_axi_gmem_cout_BREADY(m_axi_gmem_cout_BREADY),
    .m_axi_gmem_cout_BRESP(m_axi_gmem_cout_BRESP),
    .m_axi_gmem_cout_BID(m_axi_gmem_cout_BID),
    .m_axi_gmem_cout_BUSER(m_axi_gmem_cout_BUSER),
    .ap_clk(ap_clk),
    .ap_start_Boundary_X4Y12_To_X6Y12(ap_start_Boundary_X4Y12_To_X6Y12_in),
    .ap_rst_n_Boundary_X4Y12_To_X6Y12(ap_rst_n_Boundary_X4Y12_To_X6Y12_in),
    .ap_done_Boundary_X4Y12_To_X6Y12(ap_done_Boundary_X4Y12_To_X6Y12_out),
    .ap_start_Boundary_X4Y14_To_X6Y14(ap_start_Boundary_X4Y14_To_X6Y14_out),
    .ap_rst_n_Boundary_X4Y14_To_X6Y14(ap_rst_n_Boundary_X4Y14_To_X6Y14_out),
    .ap_done_Boundary_X4Y14_To_X6Y14(ap_done_Boundary_X4Y14_To_X6Y14_in)
  );


  (* keep_hierarchy = "yes" *) CR_X0Y0_To_CR_X1Y1_ctrl CR_X0Y0_To_CR_X1Y1_ctrl_U0 (
    .PE_wrapper260_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper260_U0_fifo_cin_out_V_V_din_pass_0_in),
    .PE_wrapper260_U0_fifo_cin_out_V_V_din_pass_1(PE_wrapper260_U0_fifo_cin_out_V_V_din_pass_1_out),
    .fifo_cin_PE_10_2_V_V_full_n_pass_0(fifo_cin_PE_10_2_V_V_full_n_pass_0_out),
    .fifo_cin_PE_10_2_V_V_full_n_pass_1(fifo_cin_PE_10_2_V_V_full_n_pass_1_in),
    .PE_wrapper260_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper260_U0_fifo_cin_out_V_V_write_pass_0_in),
    .PE_wrapper260_U0_fifo_cin_out_V_V_write_pass_1(PE_wrapper260_U0_fifo_cin_out_V_V_write_pass_1_out),
    .PE_wrapper261_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper261_U0_fifo_w_out_V_V_din_pass_0_in),
    .PE_wrapper261_U0_fifo_w_out_V_V_din_pass_1(PE_wrapper261_U0_fifo_w_out_V_V_din_pass_1_out),
    .fifo_w_PE_9_4_V_V_full_n_pass_0(fifo_w_PE_9_4_V_V_full_n_pass_0_out),
    .fifo_w_PE_9_4_V_V_full_n_pass_1(fifo_w_PE_9_4_V_V_full_n_pass_1_in),
    .PE_wrapper261_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper261_U0_fifo_w_out_V_V_write_pass_0_in),
    .PE_wrapper261_U0_fifo_w_out_V_V_write_pass_1(PE_wrapper261_U0_fifo_w_out_V_V_write_pass_1_out),
    .w_IO_L2_in144_U0_fifo_w_out_V_V_din_pass_0(w_IO_L2_in144_U0_fifo_w_out_V_V_din_pass_0_out),
    .fifo_w_w_IO_L2_in_10_V_V_full_n_pass_0(fifo_w_w_IO_L2_in_10_V_V_full_n_pass_0_in),
    .w_IO_L2_in144_U0_fifo_w_out_V_V_write_pass_0(w_IO_L2_in144_U0_fifo_w_out_V_V_write_pass_0_out),
    .PE_wrapper271_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper271_U0_fifo_cout_drain_out_V_din_pass_0_out),
    .fifo_cout_drain_PE_10_1_V_full_n_pass_0(fifo_cout_drain_PE_10_1_V_full_n_pass_0_in),
    .PE_wrapper271_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper271_U0_fifo_cout_drain_out_V_write_pass_0_out),
    .cout_drain_IO_L1_out_wrapper372_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper372_U0_fifo_cout_drain_out_V_V_din_pass_0_in),
    .fifo_cout_drain_cout_drain_IO_L1_out_0_10_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_0_10_V_V_full_n_pass_0_out),
    .cout_drain_IO_L1_out_wrapper372_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper372_U0_fifo_cout_drain_out_V_V_write_pass_0_in),
    .PE_wrapper247_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper247_U0_fifo_cout_drain_out_V_din_pass_0_out),
    .fifo_cout_drain_PE_8_1_V_full_n_pass_0(fifo_cout_drain_PE_8_1_V_full_n_pass_0_in),
    .PE_wrapper247_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper247_U0_fifo_cout_drain_out_V_write_pass_0_out),
    .PE_wrapper259_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper259_U0_fifo_cout_drain_out_V_din_pass_0_out),
    .fifo_cout_drain_PE_9_1_V_full_n_pass_0(fifo_cout_drain_PE_9_1_V_full_n_pass_0_in),
    .PE_wrapper259_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper259_U0_fifo_cout_drain_out_V_write_pass_0_out),
    .PE_wrapper234_U0_fifo_cin_out_V_V_din_pass_1(PE_wrapper234_U0_fifo_cin_out_V_V_din_pass_1_in),
    .fifo_cin_PE_8_0_V_V_full_n_pass_1(fifo_cin_PE_8_0_V_V_full_n_pass_1_out),
    .PE_wrapper234_U0_fifo_cin_out_V_V_write_pass_1(PE_wrapper234_U0_fifo_cin_out_V_V_write_pass_1_in),
    .PE_wrapper258_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper258_U0_fifo_cin_out_V_V_din_pass_0_out),
    .fifo_cin_PE_10_0_V_V_full_n_pass_0(fifo_cin_PE_10_0_V_V_full_n_pass_0_in),
    .PE_wrapper258_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper258_U0_fifo_cin_out_V_V_write_pass_0_out),
    .cout_drain_IO_L1_out_wrapper374_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper374_U0_fifo_cout_drain_out_V_V_din_pass_0_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_0_8_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_0_8_V_V_full_n_pass_0_in),
    .cout_drain_IO_L1_out_wrapper374_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper374_U0_fifo_cout_drain_out_V_V_write_pass_0_out),
    .PE_wrapper235_U0_fifo_cin_out_V_V_din_pass_1(PE_wrapper235_U0_fifo_cin_out_V_V_din_pass_1_in),
    .fifo_cin_PE_8_1_V_V_full_n_pass_1(fifo_cin_PE_8_1_V_V_full_n_pass_1_out),
    .PE_wrapper235_U0_fifo_cin_out_V_V_write_pass_1(PE_wrapper235_U0_fifo_cin_out_V_V_write_pass_1_in),
    .PE_wrapper247_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper247_U0_fifo_w_out_V_V_din_pass_0_out),
    .fifo_w_PE_8_2_V_V_full_n_pass_0(fifo_w_PE_8_2_V_V_full_n_pass_0_in),
    .PE_wrapper247_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper247_U0_fifo_w_out_V_V_write_pass_0_out),
    .w_IO_L2_in142_U0_fifo_w_out_V_V_din_pass_1(w_IO_L2_in142_U0_fifo_w_out_V_V_din_pass_1_in),
    .fifo_w_w_IO_L2_in_8_V_V_full_n_pass_1(fifo_w_w_IO_L2_in_8_V_V_full_n_pass_1_out),
    .w_IO_L2_in142_U0_fifo_w_out_V_V_write_pass_1(w_IO_L2_in142_U0_fifo_w_out_V_V_write_pass_1_in),
    .PE_wrapper271_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper271_U0_fifo_cin_out_V_V_din_pass_0_out),
    .fifo_cin_PE_11_1_V_V_full_n_pass_0(fifo_cin_PE_11_1_V_V_full_n_pass_0_in),
    .PE_wrapper271_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper271_U0_fifo_cin_out_V_V_write_pass_0_out),
    .PE_wrapper270_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper270_U0_fifo_w_out_V_V_din_pass_0_in),
    .fifo_w_PE_10_1_V_V_full_n_pass_0(fifo_w_PE_10_1_V_V_full_n_pass_0_out),
    .PE_wrapper270_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper270_U0_fifo_w_out_V_V_write_pass_0_in),
    .PE_wrapper259_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper259_U0_fifo_w_out_V_V_din_pass_0_out),
    .fifo_w_PE_9_2_V_V_full_n_pass_0(fifo_w_PE_9_2_V_V_full_n_pass_0_in),
    .PE_wrapper259_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper259_U0_fifo_w_out_V_V_write_pass_0_out),
    .PE_wrapper271_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper271_U0_fifo_w_out_V_V_din_pass_0_out),
    .fifo_w_PE_10_2_V_V_full_n_pass_0(fifo_w_PE_10_2_V_V_full_n_pass_0_in),
    .PE_wrapper271_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper271_U0_fifo_w_out_V_V_write_pass_0_out),
    .ap_clk(ap_clk),
    .ap_start_Boundary_X2Y0_To_X2Y2(ap_start_Boundary_X2Y0_To_X2Y2_in),
    .ap_rst_n_Boundary_X2Y0_To_X2Y2(ap_rst_n_Boundary_X2Y0_To_X2Y2_in),
    .ap_done_Boundary_X2Y0_To_X2Y2(ap_done_Boundary_X2Y0_To_X2Y2_out),
    .ap_start_Boundary_X0Y2_To_X2Y2(ap_start_Boundary_X0Y2_To_X2Y2_out),
    .ap_rst_n_Boundary_X0Y2_To_X2Y2(ap_rst_n_Boundary_X0Y2_To_X2Y2_out),
    .ap_done_Boundary_X0Y2_To_X2Y2(ap_done_Boundary_X0Y2_To_X2Y2_in)
  );


  (* keep_hierarchy = "yes" *) CR_X0Y2_To_CR_X1Y3_ctrl CR_X0Y2_To_CR_X1Y3_ctrl_U0 (
    .PE_wrapper234_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper234_U0_fifo_cin_out_V_V_din_pass_0_in),
    .PE_wrapper234_U0_fifo_cin_out_V_V_din_pass_1(PE_wrapper234_U0_fifo_cin_out_V_V_din_pass_1_out),
    .fifo_cin_PE_8_0_V_V_full_n_pass_0(fifo_cin_PE_8_0_V_V_full_n_pass_0_out),
    .fifo_cin_PE_8_0_V_V_full_n_pass_1(fifo_cin_PE_8_0_V_V_full_n_pass_1_in),
    .PE_wrapper234_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper234_U0_fifo_cin_out_V_V_write_pass_0_in),
    .PE_wrapper234_U0_fifo_cin_out_V_V_write_pass_1(PE_wrapper234_U0_fifo_cin_out_V_V_write_pass_1_out),
    .PE_wrapper235_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper235_U0_fifo_cin_out_V_V_din_pass_0_in),
    .PE_wrapper235_U0_fifo_cin_out_V_V_din_pass_1(PE_wrapper235_U0_fifo_cin_out_V_V_din_pass_1_out),
    .fifo_cin_PE_8_1_V_V_full_n_pass_0(fifo_cin_PE_8_1_V_V_full_n_pass_0_out),
    .fifo_cin_PE_8_1_V_V_full_n_pass_1(fifo_cin_PE_8_1_V_V_full_n_pass_1_in),
    .PE_wrapper235_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper235_U0_fifo_cin_out_V_V_write_pass_0_in),
    .PE_wrapper235_U0_fifo_cin_out_V_V_write_pass_1(PE_wrapper235_U0_fifo_cin_out_V_V_write_pass_1_out),
    .w_IO_L2_in142_U0_fifo_w_out_V_V_din_pass_0(w_IO_L2_in142_U0_fifo_w_out_V_V_din_pass_0_in),
    .w_IO_L2_in142_U0_fifo_w_out_V_V_din_pass_1(w_IO_L2_in142_U0_fifo_w_out_V_V_din_pass_1_out),
    .fifo_w_w_IO_L2_in_8_V_V_full_n_pass_0(fifo_w_w_IO_L2_in_8_V_V_full_n_pass_0_out),
    .fifo_w_w_IO_L2_in_8_V_V_full_n_pass_1(fifo_w_w_IO_L2_in_8_V_V_full_n_pass_1_in),
    .w_IO_L2_in142_U0_fifo_w_out_V_V_write_pass_0(w_IO_L2_in142_U0_fifo_w_out_V_V_write_pass_0_in),
    .w_IO_L2_in142_U0_fifo_w_out_V_V_write_pass_1(w_IO_L2_in142_U0_fifo_w_out_V_V_write_pass_1_out),
    .PE_wrapper261_U0_fifo_w_out_V_V_din_pass_1(PE_wrapper261_U0_fifo_w_out_V_V_din_pass_1_in),
    .PE_wrapper261_U0_fifo_w_out_V_V_din_pass_2(PE_wrapper261_U0_fifo_w_out_V_V_din_pass_2_out),
    .fifo_w_PE_9_4_V_V_full_n_pass_1(fifo_w_PE_9_4_V_V_full_n_pass_1_out),
    .fifo_w_PE_9_4_V_V_full_n_pass_2(fifo_w_PE_9_4_V_V_full_n_pass_2_in),
    .PE_wrapper261_U0_fifo_w_out_V_V_write_pass_1(PE_wrapper261_U0_fifo_w_out_V_V_write_pass_1_in),
    .PE_wrapper261_U0_fifo_w_out_V_V_write_pass_2(PE_wrapper261_U0_fifo_w_out_V_V_write_pass_2_out),
    .PE_wrapper237_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper237_U0_fifo_w_out_V_V_din_pass_0_in),
    .PE_wrapper237_U0_fifo_w_out_V_V_din_pass_1(PE_wrapper237_U0_fifo_w_out_V_V_din_pass_1_out),
    .fifo_w_PE_7_4_V_V_full_n_pass_0(fifo_w_PE_7_4_V_V_full_n_pass_0_out),
    .fifo_w_PE_7_4_V_V_full_n_pass_1(fifo_w_PE_7_4_V_V_full_n_pass_1_in),
    .PE_wrapper237_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper237_U0_fifo_w_out_V_V_write_pass_0_in),
    .PE_wrapper237_U0_fifo_w_out_V_V_write_pass_1(PE_wrapper237_U0_fifo_w_out_V_V_write_pass_1_out),
    .PE_wrapper260_U0_fifo_cin_out_V_V_din_pass_1(PE_wrapper260_U0_fifo_cin_out_V_V_din_pass_1_in),
    .fifo_cin_PE_10_2_V_V_full_n_pass_1(fifo_cin_PE_10_2_V_V_full_n_pass_1_out),
    .PE_wrapper260_U0_fifo_cin_out_V_V_write_pass_1(PE_wrapper260_U0_fifo_cin_out_V_V_write_pass_1_in),
    .cout_drain_IO_L1_out_wrapper402_U0_fifo_cout_drain_out_V_V_din_pass_2(cout_drain_IO_L1_out_wrapper402_U0_fifo_cout_drain_out_V_V_din_pass_2_in),
    .fifo_cout_drain_cout_drain_IO_L1_out_2_12_V_V_full_n_pass_2(fifo_cout_drain_cout_drain_IO_L1_out_2_12_V_V_full_n_pass_2_out),
    .cout_drain_IO_L1_out_wrapper402_U0_fifo_cout_drain_out_V_V_write_pass_2(cout_drain_IO_L1_out_wrapper402_U0_fifo_cout_drain_out_V_V_write_pass_2_in),
    .PE_wrapper271_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper271_U0_fifo_w_out_V_V_din_pass_0_in),
    .fifo_w_PE_10_2_V_V_full_n_pass_0(fifo_w_PE_10_2_V_V_full_n_pass_0_out),
    .PE_wrapper271_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper271_U0_fifo_w_out_V_V_write_pass_0_in),
    .cout_drain_IO_L1_out_wrapper372_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper372_U0_fifo_cout_drain_out_V_V_din_pass_0_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_0_10_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_0_10_V_V_full_n_pass_0_in),
    .cout_drain_IO_L1_out_wrapper372_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper372_U0_fifo_cout_drain_out_V_V_write_pass_0_out),
    .PE_wrapper247_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper247_U0_fifo_cout_drain_out_V_din_pass_0_in),
    .fifo_cout_drain_PE_8_1_V_full_n_pass_0(fifo_cout_drain_PE_8_1_V_full_n_pass_0_out),
    .PE_wrapper247_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper247_U0_fifo_cout_drain_out_V_write_pass_0_in),
    .PE_wrapper282_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper282_U0_fifo_cin_out_V_V_din_pass_0_out),
    .fifo_cin_PE_12_0_V_V_full_n_pass_0(fifo_cin_PE_12_0_V_V_full_n_pass_0_in),
    .PE_wrapper282_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper282_U0_fifo_cin_out_V_V_write_pass_0_out),
    .w_IO_L2_in146_U0_fifo_w_out_V_V_din_pass_0(w_IO_L2_in146_U0_fifo_w_out_V_V_din_pass_0_out),
    .fifo_w_w_IO_L2_in_12_V_V_full_n_pass_0(fifo_w_w_IO_L2_in_12_V_V_full_n_pass_0_in),
    .w_IO_L2_in146_U0_fifo_w_out_V_V_write_pass_0(w_IO_L2_in146_U0_fifo_w_out_V_V_write_pass_0_out),
    .PE_wrapper294_U0_fifo_cout_drain_out_V_din_pass_1(PE_wrapper294_U0_fifo_cout_drain_out_V_din_pass_1_in),
    .fifo_cout_drain_PE_12_0_V_full_n_pass_1(fifo_cout_drain_PE_12_0_V_full_n_pass_1_out),
    .PE_wrapper294_U0_fifo_cout_drain_out_V_write_pass_1(PE_wrapper294_U0_fifo_cout_drain_out_V_write_pass_1_in),
    .PE_wrapper271_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper271_U0_fifo_cin_out_V_V_din_pass_0_in),
    .fifo_cin_PE_11_1_V_V_full_n_pass_0(fifo_cin_PE_11_1_V_V_full_n_pass_0_out),
    .PE_wrapper271_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper271_U0_fifo_cin_out_V_V_write_pass_0_in),
    .w_IO_L2_in144_U0_fifo_w_out_V_V_din_pass_0(w_IO_L2_in144_U0_fifo_w_out_V_V_din_pass_0_in),
    .fifo_w_w_IO_L2_in_10_V_V_full_n_pass_0(fifo_w_w_IO_L2_in_10_V_V_full_n_pass_0_out),
    .w_IO_L2_in144_U0_fifo_w_out_V_V_write_pass_0(w_IO_L2_in144_U0_fifo_w_out_V_V_write_pass_0_in),
    .cout_drain_IO_L1_out_wrapper386_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper386_U0_fifo_cout_drain_out_V_V_din_pass_0_in),
    .fifo_cout_drain_cout_drain_IO_L1_out_1_12_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_1_12_V_V_full_n_pass_0_out),
    .cout_drain_IO_L1_out_wrapper386_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper386_U0_fifo_cout_drain_out_V_V_write_pass_0_in),
    .cout_drain_IO_L1_out_wrapper404_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper404_U0_fifo_cout_drain_out_V_V_din_pass_0_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_2_10_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_2_10_V_V_full_n_pass_0_in),
    .cout_drain_IO_L1_out_wrapper404_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper404_U0_fifo_cout_drain_out_V_V_write_pass_0_out),
    .PE_wrapper283_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper283_U0_fifo_cin_out_V_V_din_pass_0_out),
    .fifo_cin_PE_12_1_V_V_full_n_pass_0(fifo_cin_PE_12_1_V_V_full_n_pass_0_in),
    .PE_wrapper283_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper283_U0_fifo_cin_out_V_V_write_pass_0_out),
    .PE_wrapper258_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper258_U0_fifo_cin_out_V_V_din_pass_0_in),
    .fifo_cin_PE_10_0_V_V_full_n_pass_0(fifo_cin_PE_10_0_V_V_full_n_pass_0_out),
    .PE_wrapper258_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper258_U0_fifo_cin_out_V_V_write_pass_0_in),
    .cout_drain_IO_L1_out_wrapper369_U0_fifo_cout_drain_out_V_V_din_pass_1(cout_drain_IO_L1_out_wrapper369_U0_fifo_cout_drain_out_V_V_din_pass_1_in),
    .fifo_cout_drain_cout_drain_IO_L1_out_0_13_V_V_full_n_pass_1(fifo_cout_drain_cout_drain_IO_L1_out_0_13_V_V_full_n_pass_1_out),
    .cout_drain_IO_L1_out_wrapper369_U0_fifo_cout_drain_out_V_V_write_pass_1(cout_drain_IO_L1_out_wrapper369_U0_fifo_cout_drain_out_V_V_write_pass_1_in),
    .PE_wrapper270_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper270_U0_fifo_w_out_V_V_din_pass_0_out),
    .fifo_w_PE_10_1_V_V_full_n_pass_0(fifo_w_PE_10_1_V_V_full_n_pass_0_in),
    .PE_wrapper270_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper270_U0_fifo_w_out_V_V_write_pass_0_out),
    .PE_wrapper284_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper284_U0_fifo_w_out_V_V_din_pass_0_out),
    .fifo_w_PE_11_3_V_V_full_n_pass_0(fifo_w_PE_11_3_V_V_full_n_pass_0_in),
    .PE_wrapper284_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper284_U0_fifo_w_out_V_V_write_pass_0_out),
    .cout_drain_IO_L1_out_wrapper390_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper390_U0_fifo_cout_drain_out_V_V_din_pass_0_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_1_8_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_1_8_V_V_full_n_pass_0_in),
    .cout_drain_IO_L1_out_wrapper390_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper390_U0_fifo_cout_drain_out_V_V_write_pass_0_out),
    .PE_wrapper259_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper259_U0_fifo_cout_drain_out_V_din_pass_0_in),
    .fifo_cout_drain_PE_9_1_V_full_n_pass_0(fifo_cout_drain_PE_9_1_V_full_n_pass_0_out),
    .PE_wrapper259_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper259_U0_fifo_cout_drain_out_V_write_pass_0_in),
    .PE_wrapper272_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper272_U0_fifo_w_out_V_V_din_pass_0_out),
    .fifo_w_PE_10_3_V_V_full_n_pass_0(fifo_w_PE_10_3_V_V_full_n_pass_0_in),
    .PE_wrapper272_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper272_U0_fifo_w_out_V_V_write_pass_0_out),
    .PE_wrapper284_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper284_U0_fifo_cin_out_V_V_din_pass_0_out),
    .fifo_cin_PE_12_2_V_V_full_n_pass_0(fifo_cin_PE_12_2_V_V_full_n_pass_0_in),
    .PE_wrapper284_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper284_U0_fifo_cin_out_V_V_write_pass_0_out),
    .PE_wrapper271_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper271_U0_fifo_cout_drain_out_V_din_pass_0_in),
    .fifo_cout_drain_PE_10_1_V_full_n_pass_0(fifo_cout_drain_PE_10_1_V_full_n_pass_0_out),
    .PE_wrapper271_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper271_U0_fifo_cout_drain_out_V_write_pass_0_in),
    .ap_clk(ap_clk),
    .ap_start_Boundary_X0Y2_To_X2Y2(ap_start_Boundary_X0Y2_To_X2Y2_in),
    .ap_rst_n_Boundary_X0Y2_To_X2Y2(ap_rst_n_Boundary_X0Y2_To_X2Y2_in),
    .ap_done_Boundary_X0Y2_To_X2Y2(ap_done_Boundary_X0Y2_To_X2Y2_out),
    .ap_start_Boundary_X0Y4_To_X2Y4(ap_start_Boundary_X0Y4_To_X2Y4_out),
    .ap_rst_n_Boundary_X0Y4_To_X2Y4(ap_rst_n_Boundary_X0Y4_To_X2Y4_out),
    .ap_done_Boundary_X0Y4_To_X2Y4(ap_done_Boundary_X0Y4_To_X2Y4_in)
  );


  (* keep_hierarchy = "yes" *) CR_X2Y0_To_CR_X3Y1_ctrl CR_X2Y0_To_CR_X3Y1_ctrl_U0 (
    .PE_wrapper212_U0_fifo_cin_out_V_V_din_pass_1(PE_wrapper212_U0_fifo_cin_out_V_V_din_pass_1_in),
    .PE_wrapper212_U0_fifo_cin_out_V_V_din_pass_2(PE_wrapper212_U0_fifo_cin_out_V_V_din_pass_2_out),
    .fifo_cin_PE_6_2_V_V_full_n_pass_1(fifo_cin_PE_6_2_V_V_full_n_pass_1_out),
    .fifo_cin_PE_6_2_V_V_full_n_pass_2(fifo_cin_PE_6_2_V_V_full_n_pass_2_in),
    .PE_wrapper212_U0_fifo_cin_out_V_V_write_pass_1(PE_wrapper212_U0_fifo_cin_out_V_V_write_pass_1_in),
    .PE_wrapper212_U0_fifo_cin_out_V_V_write_pass_2(PE_wrapper212_U0_fifo_cin_out_V_V_write_pass_2_out),
    .PE_wrapper213_U0_fifo_cin_out_V_V_din_pass_1(PE_wrapper213_U0_fifo_cin_out_V_V_din_pass_1_in),
    .PE_wrapper213_U0_fifo_cin_out_V_V_din_pass_2(PE_wrapper213_U0_fifo_cin_out_V_V_din_pass_2_out),
    .fifo_cin_PE_6_3_V_V_full_n_pass_1(fifo_cin_PE_6_3_V_V_full_n_pass_1_out),
    .fifo_cin_PE_6_3_V_V_full_n_pass_2(fifo_cin_PE_6_3_V_V_full_n_pass_2_in),
    .PE_wrapper213_U0_fifo_cin_out_V_V_write_pass_1(PE_wrapper213_U0_fifo_cin_out_V_V_write_pass_1_in),
    .PE_wrapper213_U0_fifo_cin_out_V_V_write_pass_2(PE_wrapper213_U0_fifo_cin_out_V_V_write_pass_2_out),
    .cout_drain_IO_L1_out_wrapper374_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper374_U0_fifo_cout_drain_out_V_V_din_pass_0_in),
    .cout_drain_IO_L1_out_wrapper374_U0_fifo_cout_drain_out_V_V_din_pass_1(cout_drain_IO_L1_out_wrapper374_U0_fifo_cout_drain_out_V_V_din_pass_1_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_0_8_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_0_8_V_V_full_n_pass_0_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_0_8_V_V_full_n_pass_1(fifo_cout_drain_cout_drain_IO_L1_out_0_8_V_V_full_n_pass_1_in),
    .cout_drain_IO_L1_out_wrapper374_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper374_U0_fifo_cout_drain_out_V_V_write_pass_0_in),
    .cout_drain_IO_L1_out_wrapper374_U0_fifo_cout_drain_out_V_V_write_pass_1(cout_drain_IO_L1_out_wrapper374_U0_fifo_cout_drain_out_V_V_write_pass_1_out),
    .w_IO_L2_in140_U0_fifo_w_out_V_V_din_pass_2(w_IO_L2_in140_U0_fifo_w_out_V_V_din_pass_2_in),
    .fifo_w_w_IO_L2_in_6_V_V_full_n_pass_2(fifo_w_w_IO_L2_in_6_V_V_full_n_pass_2_out),
    .w_IO_L2_in140_U0_fifo_w_out_V_V_write_pass_2(w_IO_L2_in140_U0_fifo_w_out_V_V_write_pass_2_in),
    .PE_wrapper260_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper260_U0_fifo_cin_out_V_V_din_pass_0_out),
    .fifo_cin_PE_10_2_V_V_full_n_pass_0(fifo_cin_PE_10_2_V_V_full_n_pass_0_in),
    .PE_wrapper260_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper260_U0_fifo_cin_out_V_V_write_pass_0_out),
    .PE_wrapper224_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper224_U0_fifo_cin_out_V_V_din_pass_0_in),
    .fifo_cin_PE_7_2_V_V_full_n_pass_0(fifo_cin_PE_7_2_V_V_full_n_pass_0_out),
    .PE_wrapper224_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper224_U0_fifo_cin_out_V_V_write_pass_0_in),
    .PE_wrapper261_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper261_U0_fifo_w_out_V_V_din_pass_0_out),
    .fifo_w_PE_9_4_V_V_full_n_pass_0(fifo_w_PE_9_4_V_V_full_n_pass_0_in),
    .PE_wrapper261_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper261_U0_fifo_w_out_V_V_write_pass_0_out),
    .PE_wrapper235_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper235_U0_fifo_cout_drain_out_V_din_pass_0_in),
    .fifo_cout_drain_PE_7_1_V_full_n_pass_0(fifo_cout_drain_PE_7_1_V_full_n_pass_0_out),
    .PE_wrapper235_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper235_U0_fifo_cout_drain_out_V_write_pass_0_in),
    .PE_wrapper225_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper225_U0_fifo_cout_drain_out_V_din_pass_0_in),
    .fifo_cout_drain_PE_6_3_V_full_n_pass_0(fifo_cout_drain_PE_6_3_V_full_n_pass_0_out),
    .PE_wrapper225_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper225_U0_fifo_cout_drain_out_V_write_pass_0_in),
    .w_IO_L2_in141_U0_fifo_w_out_V_V_din_pass_0(w_IO_L2_in141_U0_fifo_w_out_V_V_din_pass_0_out),
    .fifo_w_w_IO_L2_in_7_V_V_full_n_pass_0(fifo_w_w_IO_L2_in_7_V_V_full_n_pass_0_in),
    .w_IO_L2_in141_U0_fifo_w_out_V_V_write_pass_0(w_IO_L2_in141_U0_fifo_w_out_V_V_write_pass_0_out),
    .PE_wrapper222_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper222_U0_fifo_cout_drain_out_V_din_pass_0_in),
    .fifo_cout_drain_PE_6_0_V_full_n_pass_0(fifo_cout_drain_PE_6_0_V_full_n_pass_0_out),
    .PE_wrapper222_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper222_U0_fifo_cout_drain_out_V_write_pass_0_in),
    .PE_wrapper247_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper247_U0_fifo_w_out_V_V_din_pass_0_in),
    .fifo_w_PE_8_2_V_V_full_n_pass_0(fifo_w_PE_8_2_V_V_full_n_pass_0_out),
    .PE_wrapper247_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper247_U0_fifo_w_out_V_V_write_pass_0_in),
    .cout_drain_IO_L1_out_wrapper424_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper424_U0_fifo_cout_drain_out_V_V_din_pass_0_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_3_6_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_3_6_V_V_full_n_pass_0_in),
    .cout_drain_IO_L1_out_wrapper424_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper424_U0_fifo_cout_drain_out_V_V_write_pass_0_out),
    .PE_wrapper211_U0_fifo_cin_out_V_V_din_pass_1(PE_wrapper211_U0_fifo_cin_out_V_V_din_pass_1_in),
    .fifo_cin_PE_6_1_V_V_full_n_pass_1(fifo_cin_PE_6_1_V_V_full_n_pass_1_out),
    .PE_wrapper211_U0_fifo_cin_out_V_V_write_pass_1(PE_wrapper211_U0_fifo_cin_out_V_V_write_pass_1_in),
    .cout_drain_IO_L1_out_wrapper421_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper421_U0_fifo_cout_drain_out_V_V_din_pass_0_in),
    .fifo_cout_drain_cout_drain_IO_L1_out_3_9_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_3_9_V_V_full_n_pass_0_out),
    .cout_drain_IO_L1_out_wrapper421_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper421_U0_fifo_cout_drain_out_V_V_write_pass_0_in),
    .w_IO_L2_in141_U0_fifo_w_local_out_V_V_din_pass_0(w_IO_L2_in141_U0_fifo_w_local_out_V_V_din_pass_0_out),
    .fifo_w_PE_6_0_V_V_full_n_pass_0(fifo_w_PE_6_0_V_V_full_n_pass_0_in),
    .w_IO_L2_in141_U0_fifo_w_local_out_V_V_write_pass_0(w_IO_L2_in141_U0_fifo_w_local_out_V_V_write_pass_0_out),
    .PE_wrapper261_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper261_U0_fifo_cout_drain_out_V_din_pass_0_out),
    .fifo_cout_drain_PE_9_3_V_full_n_pass_0(fifo_cout_drain_PE_9_3_V_full_n_pass_0_in),
    .PE_wrapper261_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper261_U0_fifo_cout_drain_out_V_write_pass_0_out),
    .PE_wrapper222_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper222_U0_fifo_w_out_V_V_din_pass_0_in),
    .fifo_w_PE_6_1_V_V_full_n_pass_0(fifo_w_PE_6_1_V_V_full_n_pass_0_out),
    .PE_wrapper222_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper222_U0_fifo_w_out_V_V_write_pass_0_in),
    .cout_drain_IO_L1_out_wrapper376_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper376_U0_fifo_cout_drain_out_V_V_din_pass_0_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_0_6_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_0_6_V_V_full_n_pass_0_in),
    .cout_drain_IO_L1_out_wrapper376_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper376_U0_fifo_cout_drain_out_V_V_write_pass_0_out),
    .PE_wrapper236_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper236_U0_fifo_w_out_V_V_din_pass_0_out),
    .fifo_w_PE_7_3_V_V_full_n_pass_0(fifo_w_PE_7_3_V_V_full_n_pass_0_in),
    .PE_wrapper236_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper236_U0_fifo_w_out_V_V_write_pass_0_out),
    .PE_wrapper223_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper223_U0_fifo_cin_out_V_V_din_pass_0_out),
    .fifo_cin_PE_7_1_V_V_full_n_pass_0(fifo_cin_PE_7_1_V_V_full_n_pass_0_in),
    .PE_wrapper223_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper223_U0_fifo_cin_out_V_V_write_pass_0_out),
    .cout_drain_IO_L1_out_wrapper404_U0_fifo_cout_drain_out_V_V_din_pass_1(cout_drain_IO_L1_out_wrapper404_U0_fifo_cout_drain_out_V_V_din_pass_1_in),
    .fifo_cout_drain_cout_drain_IO_L1_out_2_10_V_V_full_n_pass_1(fifo_cout_drain_cout_drain_IO_L1_out_2_10_V_V_full_n_pass_1_out),
    .cout_drain_IO_L1_out_wrapper404_U0_fifo_cout_drain_out_V_V_write_pass_1(cout_drain_IO_L1_out_wrapper404_U0_fifo_cout_drain_out_V_V_write_pass_1_in),
    .PE_wrapper249_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper249_U0_fifo_w_out_V_V_din_pass_0_out),
    .fifo_w_PE_8_4_V_V_full_n_pass_0(fifo_w_PE_8_4_V_V_full_n_pass_0_in),
    .PE_wrapper249_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper249_U0_fifo_w_out_V_V_write_pass_0_out),
    .PE_wrapper223_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper223_U0_fifo_w_out_V_V_din_pass_0_out),
    .fifo_w_PE_6_2_V_V_full_n_pass_0(fifo_w_PE_6_2_V_V_full_n_pass_0_in),
    .PE_wrapper223_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper223_U0_fifo_w_out_V_V_write_pass_0_out),
    .PE_wrapper259_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper259_U0_fifo_w_out_V_V_din_pass_0_in),
    .fifo_w_PE_9_2_V_V_full_n_pass_0(fifo_w_PE_9_2_V_V_full_n_pass_0_out),
    .PE_wrapper259_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper259_U0_fifo_w_out_V_V_write_pass_0_in),
    .cout_drain_IO_L1_out_wrapper390_U0_fifo_cout_drain_out_V_V_din_pass_1(cout_drain_IO_L1_out_wrapper390_U0_fifo_cout_drain_out_V_V_din_pass_1_in),
    .fifo_cout_drain_cout_drain_IO_L1_out_1_8_V_V_full_n_pass_1(fifo_cout_drain_cout_drain_IO_L1_out_1_8_V_V_full_n_pass_1_out),
    .cout_drain_IO_L1_out_wrapper390_U0_fifo_cout_drain_out_V_V_write_pass_1(cout_drain_IO_L1_out_wrapper390_U0_fifo_cout_drain_out_V_V_write_pass_1_in),
    .PE_wrapper237_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper237_U0_fifo_cin_out_V_V_din_pass_0_in),
    .fifo_cin_PE_8_3_V_V_full_n_pass_0(fifo_cin_PE_8_3_V_V_full_n_pass_0_out),
    .PE_wrapper237_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper237_U0_fifo_cin_out_V_V_write_pass_0_in),
    .cout_drain_IO_L1_out_wrapper408_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper408_U0_fifo_cout_drain_out_V_V_din_pass_0_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_2_6_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_2_6_V_V_full_n_pass_0_in),
    .cout_drain_IO_L1_out_wrapper408_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper408_U0_fifo_cout_drain_out_V_V_write_pass_0_out),
    .PE_wrapper224_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper224_U0_fifo_cout_drain_out_V_din_pass_0_in),
    .fifo_cout_drain_PE_6_2_V_full_n_pass_0(fifo_cout_drain_PE_6_2_V_full_n_pass_0_out),
    .PE_wrapper224_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper224_U0_fifo_cout_drain_out_V_write_pass_0_in),
    .PE_wrapper235_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper235_U0_fifo_w_out_V_V_din_pass_0_in),
    .fifo_w_PE_7_2_V_V_full_n_pass_0(fifo_w_PE_7_2_V_V_full_n_pass_0_out),
    .PE_wrapper235_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper235_U0_fifo_w_out_V_V_write_pass_0_in),
    .PE_wrapper261_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper261_U0_fifo_cin_out_V_V_din_pass_0_out),
    .fifo_cin_PE_10_3_V_V_full_n_pass_0(fifo_cin_PE_10_3_V_V_full_n_pass_0_in),
    .PE_wrapper261_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper261_U0_fifo_cin_out_V_V_write_pass_0_out),
    .cout_drain_IO_L1_out_wrapper375_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper375_U0_fifo_cout_drain_out_V_V_din_pass_0_in),
    .fifo_cout_drain_cout_drain_IO_L1_out_0_7_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_0_7_V_V_full_n_pass_0_out),
    .cout_drain_IO_L1_out_wrapper375_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper375_U0_fifo_cout_drain_out_V_V_write_pass_0_in),
    .cout_drain_IO_L1_out_wrapper392_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper392_U0_fifo_cout_drain_out_V_V_din_pass_0_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_1_6_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_1_6_V_V_full_n_pass_0_in),
    .cout_drain_IO_L1_out_wrapper392_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper392_U0_fifo_cout_drain_out_V_V_write_pass_0_out),
    .PE_wrapper237_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper237_U0_fifo_cout_drain_out_V_din_pass_0_in),
    .fifo_cout_drain_PE_7_3_V_full_n_pass_0(fifo_cout_drain_PE_7_3_V_full_n_pass_0_out),
    .PE_wrapper237_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper237_U0_fifo_cout_drain_out_V_write_pass_0_in),
    .ap_clk(ap_clk),
    .ap_start_Boundary_X4Y0_To_X4Y2(ap_start_Boundary_X4Y0_To_X4Y2_in),
    .ap_rst_n_Boundary_X4Y0_To_X4Y2(ap_rst_n_Boundary_X4Y0_To_X4Y2_in),
    .ap_done_Boundary_X4Y0_To_X4Y2(ap_done_Boundary_X4Y0_To_X4Y2_out),
    .ap_start_Boundary_X2Y2_To_X4Y2(ap_start_Boundary_X2Y2_To_X4Y2_out),
    .ap_rst_n_Boundary_X2Y2_To_X4Y2(ap_rst_n_Boundary_X2Y2_To_X4Y2_out),
    .ap_done_Boundary_X2Y2_To_X4Y2(ap_done_Boundary_X2Y2_To_X4Y2_in),
    .ap_start_Boundary_X2Y0_To_X2Y2(ap_start_Boundary_X2Y0_To_X2Y2_out),
    .ap_rst_n_Boundary_X2Y0_To_X2Y2(ap_rst_n_Boundary_X2Y0_To_X2Y2_out),
    .ap_done_Boundary_X2Y0_To_X2Y2(ap_done_Boundary_X2Y0_To_X2Y2_in)
  );


  (* keep_hierarchy = "yes" *) CR_X2Y2_To_CR_X3Y3_ctrl CR_X2Y2_To_CR_X3Y3_ctrl_U0 (
    .w_IO_L2_in140_U0_fifo_w_out_V_V_din_pass_1(w_IO_L2_in140_U0_fifo_w_out_V_V_din_pass_1_in),
    .w_IO_L2_in140_U0_fifo_w_out_V_V_din_pass_2(w_IO_L2_in140_U0_fifo_w_out_V_V_din_pass_2_out),
    .fifo_w_w_IO_L2_in_6_V_V_full_n_pass_1(fifo_w_w_IO_L2_in_6_V_V_full_n_pass_1_out),
    .fifo_w_w_IO_L2_in_6_V_V_full_n_pass_2(fifo_w_w_IO_L2_in_6_V_V_full_n_pass_2_in),
    .w_IO_L2_in140_U0_fifo_w_out_V_V_write_pass_1(w_IO_L2_in140_U0_fifo_w_out_V_V_write_pass_1_in),
    .w_IO_L2_in140_U0_fifo_w_out_V_V_write_pass_2(w_IO_L2_in140_U0_fifo_w_out_V_V_write_pass_2_out),
    .cout_drain_IO_L1_out_wrapper404_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper404_U0_fifo_cout_drain_out_V_V_din_pass_0_in),
    .cout_drain_IO_L1_out_wrapper404_U0_fifo_cout_drain_out_V_V_din_pass_1(cout_drain_IO_L1_out_wrapper404_U0_fifo_cout_drain_out_V_V_din_pass_1_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_2_10_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_2_10_V_V_full_n_pass_0_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_2_10_V_V_full_n_pass_1(fifo_cout_drain_cout_drain_IO_L1_out_2_10_V_V_full_n_pass_1_in),
    .cout_drain_IO_L1_out_wrapper404_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper404_U0_fifo_cout_drain_out_V_V_write_pass_0_in),
    .cout_drain_IO_L1_out_wrapper404_U0_fifo_cout_drain_out_V_V_write_pass_1(cout_drain_IO_L1_out_wrapper404_U0_fifo_cout_drain_out_V_V_write_pass_1_out),
    .cout_drain_IO_L1_out_wrapper390_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper390_U0_fifo_cout_drain_out_V_V_din_pass_0_in),
    .cout_drain_IO_L1_out_wrapper390_U0_fifo_cout_drain_out_V_V_din_pass_1(cout_drain_IO_L1_out_wrapper390_U0_fifo_cout_drain_out_V_V_din_pass_1_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_1_8_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_1_8_V_V_full_n_pass_0_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_1_8_V_V_full_n_pass_1(fifo_cout_drain_cout_drain_IO_L1_out_1_8_V_V_full_n_pass_1_in),
    .cout_drain_IO_L1_out_wrapper390_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper390_U0_fifo_cout_drain_out_V_V_write_pass_0_in),
    .cout_drain_IO_L1_out_wrapper390_U0_fifo_cout_drain_out_V_V_write_pass_1(cout_drain_IO_L1_out_wrapper390_U0_fifo_cout_drain_out_V_V_write_pass_1_out),
    .PE_wrapper249_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper249_U0_fifo_w_out_V_V_din_pass_0_in),
    .PE_wrapper249_U0_fifo_w_out_V_V_din_pass_1(PE_wrapper249_U0_fifo_w_out_V_V_din_pass_1_out),
    .fifo_w_PE_8_4_V_V_full_n_pass_0(fifo_w_PE_8_4_V_V_full_n_pass_0_out),
    .fifo_w_PE_8_4_V_V_full_n_pass_1(fifo_w_PE_8_4_V_V_full_n_pass_1_in),
    .PE_wrapper249_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper249_U0_fifo_w_out_V_V_write_pass_0_in),
    .PE_wrapper249_U0_fifo_w_out_V_V_write_pass_1(PE_wrapper249_U0_fifo_w_out_V_V_write_pass_1_out),
    .PE_wrapper272_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper272_U0_fifo_w_out_V_V_din_pass_0_in),
    .PE_wrapper272_U0_fifo_w_out_V_V_din_pass_1(PE_wrapper272_U0_fifo_w_out_V_V_din_pass_1_out),
    .fifo_w_PE_10_3_V_V_full_n_pass_0(fifo_w_PE_10_3_V_V_full_n_pass_0_out),
    .fifo_w_PE_10_3_V_V_full_n_pass_1(fifo_w_PE_10_3_V_V_full_n_pass_1_in),
    .PE_wrapper272_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper272_U0_fifo_w_out_V_V_write_pass_0_in),
    .PE_wrapper272_U0_fifo_w_out_V_V_write_pass_1(PE_wrapper272_U0_fifo_w_out_V_V_write_pass_1_out),
    .PE_wrapper261_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper261_U0_fifo_cin_out_V_V_din_pass_0_in),
    .PE_wrapper261_U0_fifo_cin_out_V_V_din_pass_1(PE_wrapper261_U0_fifo_cin_out_V_V_din_pass_1_out),
    .fifo_cin_PE_10_3_V_V_full_n_pass_0(fifo_cin_PE_10_3_V_V_full_n_pass_0_out),
    .fifo_cin_PE_10_3_V_V_full_n_pass_1(fifo_cin_PE_10_3_V_V_full_n_pass_1_in),
    .PE_wrapper261_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper261_U0_fifo_cin_out_V_V_write_pass_0_in),
    .PE_wrapper261_U0_fifo_cin_out_V_V_write_pass_1(PE_wrapper261_U0_fifo_cin_out_V_V_write_pass_1_out),
    .PE_wrapper224_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper224_U0_fifo_cin_out_V_V_din_pass_0_out),
    .fifo_cin_PE_7_2_V_V_full_n_pass_0(fifo_cin_PE_7_2_V_V_full_n_pass_0_in),
    .PE_wrapper224_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper224_U0_fifo_cin_out_V_V_write_pass_0_out),
    .PE_wrapper235_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper235_U0_fifo_cout_drain_out_V_din_pass_0_out),
    .fifo_cout_drain_PE_7_1_V_full_n_pass_0(fifo_cout_drain_PE_7_1_V_full_n_pass_0_in),
    .PE_wrapper235_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper235_U0_fifo_cout_drain_out_V_write_pass_0_out),
    .PE_wrapper225_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper225_U0_fifo_cout_drain_out_V_din_pass_0_out),
    .fifo_cout_drain_PE_6_3_V_full_n_pass_0(fifo_cout_drain_PE_6_3_V_full_n_pass_0_in),
    .PE_wrapper225_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper225_U0_fifo_cout_drain_out_V_write_pass_0_out),
    .w_IO_L2_in141_U0_fifo_w_out_V_V_din_pass_0(w_IO_L2_in141_U0_fifo_w_out_V_V_din_pass_0_in),
    .fifo_w_w_IO_L2_in_7_V_V_full_n_pass_0(fifo_w_w_IO_L2_in_7_V_V_full_n_pass_0_out),
    .w_IO_L2_in141_U0_fifo_w_out_V_V_write_pass_0(w_IO_L2_in141_U0_fifo_w_out_V_V_write_pass_0_in),
    .PE_wrapper235_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper235_U0_fifo_cin_out_V_V_din_pass_0_out),
    .fifo_cin_PE_8_1_V_V_full_n_pass_0(fifo_cin_PE_8_1_V_V_full_n_pass_0_in),
    .PE_wrapper235_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper235_U0_fifo_cin_out_V_V_write_pass_0_out),
    .PE_wrapper222_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper222_U0_fifo_cout_drain_out_V_din_pass_0_out),
    .fifo_cout_drain_PE_6_0_V_full_n_pass_0(fifo_cout_drain_PE_6_0_V_full_n_pass_0_in),
    .PE_wrapper222_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper222_U0_fifo_cout_drain_out_V_write_pass_0_out),
    .PE_wrapper212_U0_fifo_cin_out_V_V_din_pass_2(PE_wrapper212_U0_fifo_cin_out_V_V_din_pass_2_in),
    .fifo_cin_PE_6_2_V_V_full_n_pass_2(fifo_cin_PE_6_2_V_V_full_n_pass_2_out),
    .PE_wrapper212_U0_fifo_cin_out_V_V_write_pass_2(PE_wrapper212_U0_fifo_cin_out_V_V_write_pass_2_in),
    .PE_wrapper225_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper225_U0_fifo_w_out_V_V_din_pass_0_out),
    .fifo_w_PE_6_4_V_V_full_n_pass_0(fifo_w_PE_6_4_V_V_full_n_pass_0_in),
    .PE_wrapper225_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper225_U0_fifo_w_out_V_V_write_pass_0_out),
    .cout_drain_IO_L1_out_wrapper421_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper421_U0_fifo_cout_drain_out_V_V_din_pass_0_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_3_9_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_3_9_V_V_full_n_pass_0_in),
    .cout_drain_IO_L1_out_wrapper421_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper421_U0_fifo_cout_drain_out_V_V_write_pass_0_out),
    .w_IO_L2_in141_U0_fifo_w_local_out_V_V_din_pass_0(w_IO_L2_in141_U0_fifo_w_local_out_V_V_din_pass_0_in),
    .fifo_w_PE_6_0_V_V_full_n_pass_0(fifo_w_PE_6_0_V_V_full_n_pass_0_out),
    .w_IO_L2_in141_U0_fifo_w_local_out_V_V_write_pass_0(w_IO_L2_in141_U0_fifo_w_local_out_V_V_write_pass_0_in),
    .cout_drain_IO_L1_out_wrapper375_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper375_U0_fifo_cout_drain_out_V_V_din_pass_0_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_0_7_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_0_7_V_V_full_n_pass_0_in),
    .cout_drain_IO_L1_out_wrapper375_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper375_U0_fifo_cout_drain_out_V_V_write_pass_0_out),
    .PE_wrapper261_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper261_U0_fifo_cout_drain_out_V_din_pass_0_in),
    .fifo_cout_drain_PE_9_3_V_full_n_pass_0(fifo_cout_drain_PE_9_3_V_full_n_pass_0_out),
    .PE_wrapper261_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper261_U0_fifo_cout_drain_out_V_write_pass_0_in),
    .PE_wrapper213_U0_fifo_cin_out_V_V_din_pass_2(PE_wrapper213_U0_fifo_cin_out_V_V_din_pass_2_in),
    .fifo_cin_PE_6_3_V_V_full_n_pass_2(fifo_cin_PE_6_3_V_V_full_n_pass_2_out),
    .PE_wrapper213_U0_fifo_cin_out_V_V_write_pass_2(PE_wrapper213_U0_fifo_cin_out_V_V_write_pass_2_in),
    .PE_wrapper222_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper222_U0_fifo_w_out_V_V_din_pass_0_out),
    .fifo_w_PE_6_1_V_V_full_n_pass_0(fifo_w_PE_6_1_V_V_full_n_pass_0_in),
    .PE_wrapper222_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper222_U0_fifo_w_out_V_V_write_pass_0_out),
    .PE_wrapper237_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper237_U0_fifo_w_out_V_V_din_pass_0_out),
    .fifo_w_PE_7_4_V_V_full_n_pass_0(fifo_w_PE_7_4_V_V_full_n_pass_0_in),
    .PE_wrapper237_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper237_U0_fifo_w_out_V_V_write_pass_0_out),
    .PE_wrapper236_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper236_U0_fifo_w_out_V_V_din_pass_0_in),
    .fifo_w_PE_7_3_V_V_full_n_pass_0(fifo_w_PE_7_3_V_V_full_n_pass_0_out),
    .PE_wrapper236_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper236_U0_fifo_w_out_V_V_write_pass_0_in),
    .PE_wrapper223_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper223_U0_fifo_cin_out_V_V_din_pass_0_in),
    .fifo_cin_PE_7_1_V_V_full_n_pass_0(fifo_cin_PE_7_1_V_V_full_n_pass_0_out),
    .PE_wrapper223_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper223_U0_fifo_cin_out_V_V_write_pass_0_in),
    .cout_drain_IO_L1_out_wrapper374_U0_fifo_cout_drain_out_V_V_din_pass_1(cout_drain_IO_L1_out_wrapper374_U0_fifo_cout_drain_out_V_V_din_pass_1_in),
    .fifo_cout_drain_cout_drain_IO_L1_out_0_8_V_V_full_n_pass_1(fifo_cout_drain_cout_drain_IO_L1_out_0_8_V_V_full_n_pass_1_out),
    .cout_drain_IO_L1_out_wrapper374_U0_fifo_cout_drain_out_V_V_write_pass_1(cout_drain_IO_L1_out_wrapper374_U0_fifo_cout_drain_out_V_V_write_pass_1_in),
    .PE_wrapper223_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper223_U0_fifo_w_out_V_V_din_pass_0_in),
    .fifo_w_PE_6_2_V_V_full_n_pass_0(fifo_w_PE_6_2_V_V_full_n_pass_0_out),
    .PE_wrapper223_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper223_U0_fifo_w_out_V_V_write_pass_0_in),
    .cout_drain_IO_L1_out_wrapper420_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper420_U0_fifo_cout_drain_out_V_V_din_pass_0_in),
    .fifo_cout_drain_cout_drain_IO_L1_out_3_10_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_3_10_V_V_full_n_pass_0_out),
    .cout_drain_IO_L1_out_wrapper420_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper420_U0_fifo_cout_drain_out_V_V_write_pass_0_in),
    .PE_wrapper234_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper234_U0_fifo_cin_out_V_V_din_pass_0_out),
    .fifo_cin_PE_8_0_V_V_full_n_pass_0(fifo_cin_PE_8_0_V_V_full_n_pass_0_in),
    .PE_wrapper234_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper234_U0_fifo_cin_out_V_V_write_pass_0_out),
    .PE_wrapper237_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper237_U0_fifo_cin_out_V_V_din_pass_0_out),
    .fifo_cin_PE_8_3_V_V_full_n_pass_0(fifo_cin_PE_8_3_V_V_full_n_pass_0_in),
    .PE_wrapper237_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper237_U0_fifo_cin_out_V_V_write_pass_0_out),
    .PE_wrapper235_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper235_U0_fifo_w_out_V_V_din_pass_0_out),
    .fifo_w_PE_7_2_V_V_full_n_pass_0(fifo_w_PE_7_2_V_V_full_n_pass_0_in),
    .PE_wrapper235_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper235_U0_fifo_w_out_V_V_write_pass_0_out),
    .w_IO_L2_in142_U0_fifo_w_out_V_V_din_pass_0(w_IO_L2_in142_U0_fifo_w_out_V_V_din_pass_0_out),
    .fifo_w_w_IO_L2_in_8_V_V_full_n_pass_0(fifo_w_w_IO_L2_in_8_V_V_full_n_pass_0_in),
    .w_IO_L2_in142_U0_fifo_w_out_V_V_write_pass_0(w_IO_L2_in142_U0_fifo_w_out_V_V_write_pass_0_out),
    .PE_wrapper224_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper224_U0_fifo_cout_drain_out_V_din_pass_0_out),
    .fifo_cout_drain_PE_6_2_V_full_n_pass_0(fifo_cout_drain_PE_6_2_V_full_n_pass_0_in),
    .PE_wrapper224_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper224_U0_fifo_cout_drain_out_V_write_pass_0_out),
    .PE_wrapper210_U0_fifo_cin_out_V_V_din_pass_1(PE_wrapper210_U0_fifo_cin_out_V_V_din_pass_1_in),
    .fifo_cin_PE_6_0_V_V_full_n_pass_1(fifo_cin_PE_6_0_V_V_full_n_pass_1_out),
    .PE_wrapper210_U0_fifo_cin_out_V_V_write_pass_1(PE_wrapper210_U0_fifo_cin_out_V_V_write_pass_1_in),
    .PE_wrapper237_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper237_U0_fifo_cout_drain_out_V_din_pass_0_out),
    .fifo_cout_drain_PE_7_3_V_full_n_pass_0(fifo_cout_drain_PE_7_3_V_full_n_pass_0_in),
    .PE_wrapper237_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper237_U0_fifo_cout_drain_out_V_write_pass_0_out),
    .ap_clk(ap_clk),
    .ap_start_Boundary_X2Y2_To_X4Y2(ap_start_Boundary_X2Y2_To_X4Y2_in),
    .ap_rst_n_Boundary_X2Y2_To_X4Y2(ap_rst_n_Boundary_X2Y2_To_X4Y2_in),
    .ap_done_Boundary_X2Y2_To_X4Y2(ap_done_Boundary_X2Y2_To_X4Y2_out),
    .ap_start_Boundary_X2Y4_To_X4Y4(ap_start_Boundary_X2Y4_To_X4Y4_out),
    .ap_rst_n_Boundary_X2Y4_To_X4Y4(ap_rst_n_Boundary_X2Y4_To_X4Y4_out),
    .ap_done_Boundary_X2Y4_To_X4Y4(ap_done_Boundary_X2Y4_To_X4Y4_in)
  );


  (* keep_hierarchy = "yes" *) CR_X0Y4_To_CR_X1Y5_ctrl CR_X0Y4_To_CR_X1Y5_ctrl_U0 (
    .cout_drain_IO_L1_out_wrapper402_U0_fifo_cout_drain_out_V_V_din_pass_1(cout_drain_IO_L1_out_wrapper402_U0_fifo_cout_drain_out_V_V_din_pass_1_in),
    .cout_drain_IO_L1_out_wrapper402_U0_fifo_cout_drain_out_V_V_din_pass_2(cout_drain_IO_L1_out_wrapper402_U0_fifo_cout_drain_out_V_V_din_pass_2_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_2_12_V_V_full_n_pass_1(fifo_cout_drain_cout_drain_IO_L1_out_2_12_V_V_full_n_pass_1_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_2_12_V_V_full_n_pass_2(fifo_cout_drain_cout_drain_IO_L1_out_2_12_V_V_full_n_pass_2_in),
    .cout_drain_IO_L1_out_wrapper402_U0_fifo_cout_drain_out_V_V_write_pass_1(cout_drain_IO_L1_out_wrapper402_U0_fifo_cout_drain_out_V_V_write_pass_1_in),
    .cout_drain_IO_L1_out_wrapper402_U0_fifo_cout_drain_out_V_V_write_pass_2(cout_drain_IO_L1_out_wrapper402_U0_fifo_cout_drain_out_V_V_write_pass_2_out),
    .PE_wrapper294_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper294_U0_fifo_cout_drain_out_V_din_pass_0_in),
    .PE_wrapper294_U0_fifo_cout_drain_out_V_din_pass_1(PE_wrapper294_U0_fifo_cout_drain_out_V_din_pass_1_out),
    .fifo_cout_drain_PE_12_0_V_full_n_pass_0(fifo_cout_drain_PE_12_0_V_full_n_pass_0_out),
    .fifo_cout_drain_PE_12_0_V_full_n_pass_1(fifo_cout_drain_PE_12_0_V_full_n_pass_1_in),
    .PE_wrapper294_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper294_U0_fifo_cout_drain_out_V_write_pass_0_in),
    .PE_wrapper294_U0_fifo_cout_drain_out_V_write_pass_1(PE_wrapper294_U0_fifo_cout_drain_out_V_write_pass_1_out),
    .cout_drain_IO_L1_out_wrapper369_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper369_U0_fifo_cout_drain_out_V_V_din_pass_0_in),
    .cout_drain_IO_L1_out_wrapper369_U0_fifo_cout_drain_out_V_V_din_pass_1(cout_drain_IO_L1_out_wrapper369_U0_fifo_cout_drain_out_V_V_din_pass_1_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_0_13_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_0_13_V_V_full_n_pass_0_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_0_13_V_V_full_n_pass_1(fifo_cout_drain_cout_drain_IO_L1_out_0_13_V_V_full_n_pass_1_in),
    .cout_drain_IO_L1_out_wrapper369_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper369_U0_fifo_cout_drain_out_V_V_write_pass_0_in),
    .cout_drain_IO_L1_out_wrapper369_U0_fifo_cout_drain_out_V_V_write_pass_1(cout_drain_IO_L1_out_wrapper369_U0_fifo_cout_drain_out_V_V_write_pass_1_out),
    .PE_wrapper298_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper298_U0_fifo_cin_out_V_V_din_pass_0_in),
    .PE_wrapper298_U0_fifo_cin_out_V_V_din_pass_1(PE_wrapper298_U0_fifo_cin_out_V_V_din_pass_1_out),
    .fifo_cin_PE_13_4_V_V_full_n_pass_0(fifo_cin_PE_13_4_V_V_full_n_pass_0_out),
    .fifo_cin_PE_13_4_V_V_full_n_pass_1(fifo_cin_PE_13_4_V_V_full_n_pass_1_in),
    .PE_wrapper298_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper298_U0_fifo_cin_out_V_V_write_pass_0_in),
    .PE_wrapper298_U0_fifo_cin_out_V_V_write_pass_1(PE_wrapper298_U0_fifo_cin_out_V_V_write_pass_1_out),
    .PE_wrapper250_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper250_U0_fifo_cout_drain_out_V_din_pass_0_in),
    .PE_wrapper250_U0_fifo_cout_drain_out_V_din_pass_1(PE_wrapper250_U0_fifo_cout_drain_out_V_din_pass_1_out),
    .fifo_cout_drain_PE_8_4_V_full_n_pass_0(fifo_cout_drain_PE_8_4_V_full_n_pass_0_out),
    .fifo_cout_drain_PE_8_4_V_full_n_pass_1(fifo_cout_drain_PE_8_4_V_full_n_pass_1_in),
    .PE_wrapper250_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper250_U0_fifo_cout_drain_out_V_write_pass_0_in),
    .PE_wrapper250_U0_fifo_cout_drain_out_V_write_pass_1(PE_wrapper250_U0_fifo_cout_drain_out_V_write_pass_1_out),
    .PE_wrapper282_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper282_U0_fifo_cin_out_V_V_din_pass_0_in),
    .PE_wrapper282_U0_fifo_cin_out_V_V_din_pass_1(PE_wrapper282_U0_fifo_cin_out_V_V_din_pass_1_out),
    .fifo_cin_PE_12_0_V_V_full_n_pass_0(fifo_cin_PE_12_0_V_V_full_n_pass_0_out),
    .fifo_cin_PE_12_0_V_V_full_n_pass_1(fifo_cin_PE_12_0_V_V_full_n_pass_1_in),
    .PE_wrapper282_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper282_U0_fifo_cin_out_V_V_write_pass_0_in),
    .PE_wrapper282_U0_fifo_cin_out_V_V_write_pass_1(PE_wrapper282_U0_fifo_cin_out_V_V_write_pass_1_out),
    .PE_wrapper237_U0_fifo_w_out_V_V_din_pass_1(PE_wrapper237_U0_fifo_w_out_V_V_din_pass_1_in),
    .PE_wrapper237_U0_fifo_w_out_V_V_din_pass_2(PE_wrapper237_U0_fifo_w_out_V_V_din_pass_2_out),
    .fifo_w_PE_7_4_V_V_full_n_pass_1(fifo_w_PE_7_4_V_V_full_n_pass_1_out),
    .fifo_w_PE_7_4_V_V_full_n_pass_2(fifo_w_PE_7_4_V_V_full_n_pass_2_in),
    .PE_wrapper237_U0_fifo_w_out_V_V_write_pass_1(PE_wrapper237_U0_fifo_w_out_V_V_write_pass_1_in),
    .PE_wrapper237_U0_fifo_w_out_V_V_write_pass_2(PE_wrapper237_U0_fifo_w_out_V_V_write_pass_2_out),
    .PE_wrapper283_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper283_U0_fifo_cin_out_V_V_din_pass_0_in),
    .PE_wrapper283_U0_fifo_cin_out_V_V_din_pass_1(PE_wrapper283_U0_fifo_cin_out_V_V_din_pass_1_out),
    .fifo_cin_PE_12_1_V_V_full_n_pass_0(fifo_cin_PE_12_1_V_V_full_n_pass_0_out),
    .fifo_cin_PE_12_1_V_V_full_n_pass_1(fifo_cin_PE_12_1_V_V_full_n_pass_1_in),
    .PE_wrapper283_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper283_U0_fifo_cin_out_V_V_write_pass_0_in),
    .PE_wrapper283_U0_fifo_cin_out_V_V_write_pass_1(PE_wrapper283_U0_fifo_cin_out_V_V_write_pass_1_out),
    .PE_wrapper298_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper298_U0_fifo_w_out_V_V_din_pass_0_in),
    .PE_wrapper298_U0_fifo_w_out_V_V_din_pass_1(PE_wrapper298_U0_fifo_w_out_V_V_din_pass_1_out),
    .fifo_w_PE_12_5_V_V_full_n_pass_0(fifo_w_PE_12_5_V_V_full_n_pass_0_out),
    .fifo_w_PE_12_5_V_V_full_n_pass_1(fifo_w_PE_12_5_V_V_full_n_pass_1_in),
    .PE_wrapper298_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper298_U0_fifo_w_out_V_V_write_pass_0_in),
    .PE_wrapper298_U0_fifo_w_out_V_V_write_pass_1(PE_wrapper298_U0_fifo_w_out_V_V_write_pass_1_out),
    .PE_wrapper322_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper322_U0_fifo_w_out_V_V_din_pass_0_in),
    .PE_wrapper322_U0_fifo_w_out_V_V_din_pass_1(PE_wrapper322_U0_fifo_w_out_V_V_din_pass_1_out),
    .fifo_w_PE_14_5_V_V_full_n_pass_0(fifo_w_PE_14_5_V_V_full_n_pass_0_out),
    .fifo_w_PE_14_5_V_V_full_n_pass_1(fifo_w_PE_14_5_V_V_full_n_pass_1_in),
    .PE_wrapper322_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper322_U0_fifo_w_out_V_V_write_pass_0_in),
    .PE_wrapper322_U0_fifo_w_out_V_V_write_pass_1(PE_wrapper322_U0_fifo_w_out_V_V_write_pass_1_out),
    .PE_wrapper334_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper334_U0_fifo_w_out_V_V_din_pass_0_in),
    .PE_wrapper334_U0_fifo_w_out_V_V_din_pass_1(PE_wrapper334_U0_fifo_w_out_V_V_din_pass_1_out),
    .fifo_w_PE_15_5_V_V_full_n_pass_0(fifo_w_PE_15_5_V_V_full_n_pass_0_out),
    .fifo_w_PE_15_5_V_V_full_n_pass_1(fifo_w_PE_15_5_V_V_full_n_pass_1_in),
    .PE_wrapper334_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper334_U0_fifo_w_out_V_V_write_pass_0_in),
    .PE_wrapper334_U0_fifo_w_out_V_V_write_pass_1(PE_wrapper334_U0_fifo_w_out_V_V_write_pass_1_out),
    .cout_drain_IO_L1_out_wrapper385_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper385_U0_fifo_cout_drain_out_V_V_din_pass_0_in),
    .fifo_cout_drain_cout_drain_IO_L1_out_1_13_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_1_13_V_V_full_n_pass_0_out),
    .cout_drain_IO_L1_out_wrapper385_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper385_U0_fifo_cout_drain_out_V_V_write_pass_0_in),
    .PE_wrapper309_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper309_U0_fifo_cin_out_V_V_din_pass_0_out),
    .fifo_cin_PE_14_3_V_V_full_n_pass_0(fifo_cin_PE_14_3_V_V_full_n_pass_0_in),
    .PE_wrapper309_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper309_U0_fifo_cin_out_V_V_write_pass_0_out),
    .PE_wrapper261_U0_fifo_w_out_V_V_din_pass_2(PE_wrapper261_U0_fifo_w_out_V_V_din_pass_2_in),
    .fifo_w_PE_9_4_V_V_full_n_pass_2(fifo_w_PE_9_4_V_V_full_n_pass_2_out),
    .PE_wrapper261_U0_fifo_w_out_V_V_write_pass_2(PE_wrapper261_U0_fifo_w_out_V_V_write_pass_2_in),
    .PE_wrapper333_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper333_U0_fifo_w_out_V_V_din_pass_0_out),
    .fifo_w_PE_15_4_V_V_full_n_pass_0(fifo_w_PE_15_4_V_V_full_n_pass_0_in),
    .PE_wrapper333_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper333_U0_fifo_w_out_V_V_write_pass_0_out),
    .cout_drain_IO_L1_out_wrapper440_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper440_U0_fifo_cout_drain_out_V_V_din_pass_0_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_4_6_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_4_6_V_V_full_n_pass_0_in),
    .cout_drain_IO_L1_out_wrapper440_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper440_U0_fifo_cout_drain_out_V_V_write_pass_0_out),
    .PE_wrapper250_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper250_U0_fifo_cin_out_V_V_din_pass_0_in),
    .fifo_cin_PE_9_4_V_V_full_n_pass_0(fifo_cin_PE_9_4_V_V_full_n_pass_0_out),
    .PE_wrapper250_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper250_U0_fifo_cin_out_V_V_write_pass_0_in),
    .PE_wrapper286_U0_fifo_cout_drain_out_V_din_pass_1(PE_wrapper286_U0_fifo_cout_drain_out_V_din_pass_1_in),
    .fifo_cout_drain_PE_11_4_V_full_n_pass_1(fifo_cout_drain_PE_11_4_V_full_n_pass_1_out),
    .PE_wrapper286_U0_fifo_cout_drain_out_V_write_pass_1(PE_wrapper286_U0_fifo_cout_drain_out_V_write_pass_1_in),
    .cout_drain_IO_L1_out_wrapper439_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper439_U0_fifo_cout_drain_out_V_V_din_pass_0_in),
    .fifo_cout_drain_cout_drain_IO_L1_out_4_7_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_4_7_V_V_full_n_pass_0_out),
    .cout_drain_IO_L1_out_wrapper439_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper439_U0_fifo_cout_drain_out_V_V_write_pass_0_in),
    .PE_wrapper306_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper306_U0_fifo_cout_drain_out_V_din_pass_0_out),
    .fifo_cout_drain_PE_13_0_V_full_n_pass_0(fifo_cout_drain_PE_13_0_V_full_n_pass_0_in),
    .PE_wrapper306_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper306_U0_fifo_cout_drain_out_V_write_pass_0_out),
    .PE_wrapper295_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper295_U0_fifo_w_out_V_V_din_pass_0_in),
    .fifo_w_PE_12_2_V_V_full_n_pass_0(fifo_w_PE_12_2_V_V_full_n_pass_0_out),
    .PE_wrapper295_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper295_U0_fifo_w_out_V_V_write_pass_0_in),
    .PE_wrapper226_U0_fifo_cout_drain_out_V_din_pass_1(PE_wrapper226_U0_fifo_cout_drain_out_V_din_pass_1_in),
    .fifo_cout_drain_PE_6_4_V_full_n_pass_1(fifo_cout_drain_PE_6_4_V_full_n_pass_1_out),
    .PE_wrapper226_U0_fifo_cout_drain_out_V_write_pass_1(PE_wrapper226_U0_fifo_cout_drain_out_V_write_pass_1_in),
    .PE_wrapper320_U0_fifo_cin_out_V_V_din_pass_1(PE_wrapper320_U0_fifo_cin_out_V_V_din_pass_1_in),
    .fifo_cin_PE_15_2_V_V_full_n_pass_1(fifo_cin_PE_15_2_V_V_full_n_pass_1_out),
    .PE_wrapper320_U0_fifo_cin_out_V_V_write_pass_1(PE_wrapper320_U0_fifo_cin_out_V_V_write_pass_1_in),
    .PE_wrapper309_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper309_U0_fifo_w_out_V_V_din_pass_0_out),
    .fifo_w_PE_13_4_V_V_full_n_pass_0(fifo_w_PE_13_4_V_V_full_n_pass_0_in),
    .PE_wrapper309_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper309_U0_fifo_w_out_V_V_write_pass_0_out),
    .PE_wrapper331_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper331_U0_fifo_w_out_V_V_din_pass_0_in),
    .fifo_w_PE_15_2_V_V_full_n_pass_0(fifo_w_PE_15_2_V_V_full_n_pass_0_out),
    .PE_wrapper331_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper331_U0_fifo_w_out_V_V_write_pass_0_in),
    .cout_drain_IO_L1_out_wrapper418_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper418_U0_fifo_cout_drain_out_V_V_din_pass_0_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_3_12_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_3_12_V_V_full_n_pass_0_in),
    .cout_drain_IO_L1_out_wrapper418_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper418_U0_fifo_cout_drain_out_V_V_write_pass_0_out),
    .cout_drain_IO_L1_out_wrapper417_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper417_U0_fifo_cout_drain_out_V_V_din_pass_0_in),
    .fifo_cout_drain_cout_drain_IO_L1_out_3_13_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_3_13_V_V_full_n_pass_0_out),
    .cout_drain_IO_L1_out_wrapper417_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper417_U0_fifo_cout_drain_out_V_V_write_pass_0_in),
    .w_IO_L2_in147_U0_fifo_w_out_V_V_din_pass_0(w_IO_L2_in147_U0_fifo_w_out_V_V_din_pass_0_out),
    .fifo_w_w_IO_L2_in_13_V_V_full_n_pass_0(fifo_w_w_IO_L2_in_13_V_V_full_n_pass_0_in),
    .w_IO_L2_in147_U0_fifo_w_out_V_V_write_pass_0(w_IO_L2_in147_U0_fifo_w_out_V_V_write_pass_0_out),
    .w_IO_L2_in146_U0_fifo_w_out_V_V_din_pass_0(w_IO_L2_in146_U0_fifo_w_out_V_V_din_pass_0_in),
    .fifo_w_w_IO_L2_in_12_V_V_full_n_pass_0(fifo_w_w_IO_L2_in_12_V_V_full_n_pass_0_out),
    .w_IO_L2_in146_U0_fifo_w_out_V_V_write_pass_0(w_IO_L2_in146_U0_fifo_w_out_V_V_write_pass_0_in),
    .PE_wrapper297_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper297_U0_fifo_cin_out_V_V_din_pass_0_in),
    .fifo_cin_PE_13_3_V_V_full_n_pass_0(fifo_cin_PE_13_3_V_V_full_n_pass_0_out),
    .PE_wrapper297_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper297_U0_fifo_cin_out_V_V_write_pass_0_in),
    .PE_wrapper285_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper285_U0_fifo_w_out_V_V_din_pass_0_out),
    .fifo_w_PE_11_4_V_V_full_n_pass_0(fifo_w_PE_11_4_V_V_full_n_pass_0_in),
    .PE_wrapper285_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper285_U0_fifo_w_out_V_V_write_pass_0_out),
    .PE_wrapper306_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper306_U0_fifo_w_out_V_V_din_pass_0_out),
    .fifo_w_PE_13_1_V_V_full_n_pass_0(fifo_w_PE_13_1_V_V_full_n_pass_0_in),
    .PE_wrapper306_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper306_U0_fifo_w_out_V_V_write_pass_0_out),
    .PE_wrapper333_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper333_U0_fifo_cout_drain_out_V_din_pass_0_out),
    .fifo_cout_drain_PE_15_3_V_full_n_pass_0(fifo_cout_drain_PE_15_3_V_full_n_pass_0_in),
    .PE_wrapper333_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper333_U0_fifo_cout_drain_out_V_write_pass_0_out),
    .cout_drain_IO_L1_out_wrapper386_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper386_U0_fifo_cout_drain_out_V_V_din_pass_0_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_1_12_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_1_12_V_V_full_n_pass_0_in),
    .cout_drain_IO_L1_out_wrapper386_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper386_U0_fifo_cout_drain_out_V_V_write_pass_0_out),
    .PE_wrapper262_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper262_U0_fifo_w_out_V_V_din_pass_0_out),
    .fifo_w_PE_9_5_V_V_full_n_pass_0(fifo_w_PE_9_5_V_V_full_n_pass_0_in),
    .PE_wrapper262_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper262_U0_fifo_w_out_V_V_write_pass_0_out),
    .PE_wrapper306_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper306_U0_fifo_cin_out_V_V_din_pass_0_out),
    .fifo_cin_PE_14_0_V_V_full_n_pass_0(fifo_cin_PE_14_0_V_V_full_n_pass_0_in),
    .PE_wrapper306_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper306_U0_fifo_cin_out_V_V_write_pass_0_out),
    .PE_wrapper273_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper273_U0_fifo_cin_out_V_V_din_pass_0_in),
    .fifo_cin_PE_11_3_V_V_full_n_pass_0(fifo_cin_PE_11_3_V_V_full_n_pass_0_out),
    .PE_wrapper273_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper273_U0_fifo_cin_out_V_V_write_pass_0_in),
    .PE_wrapper321_U0_fifo_cin_out_V_V_din_pass_1(PE_wrapper321_U0_fifo_cin_out_V_V_din_pass_1_in),
    .fifo_cin_PE_15_3_V_V_full_n_pass_1(fifo_cin_PE_15_3_V_V_full_n_pass_1_out),
    .PE_wrapper321_U0_fifo_cin_out_V_V_write_pass_1(PE_wrapper321_U0_fifo_cin_out_V_V_write_pass_1_in),
    .PE_wrapper295_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper295_U0_fifo_cout_drain_out_V_din_pass_0_in),
    .fifo_cout_drain_PE_12_1_V_full_n_pass_0(fifo_cout_drain_PE_12_1_V_full_n_pass_0_out),
    .PE_wrapper295_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper295_U0_fifo_cout_drain_out_V_write_pass_0_in),
    .PE_wrapper285_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper285_U0_fifo_cout_drain_out_V_din_pass_0_out),
    .fifo_cout_drain_PE_11_3_V_full_n_pass_0(fifo_cout_drain_PE_11_3_V_full_n_pass_0_in),
    .PE_wrapper285_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper285_U0_fifo_cout_drain_out_V_write_pass_0_out),
    .PE_wrapper294_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper294_U0_fifo_cin_out_V_V_din_pass_0_in),
    .fifo_cin_PE_13_0_V_V_full_n_pass_0(fifo_cin_PE_13_0_V_V_full_n_pass_0_out),
    .PE_wrapper294_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper294_U0_fifo_cin_out_V_V_write_pass_0_in),
    .w_IO_L2_in147_U0_fifo_w_local_out_V_V_din_pass_0(w_IO_L2_in147_U0_fifo_w_local_out_V_V_din_pass_0_out),
    .fifo_w_PE_12_0_V_V_full_n_pass_0(fifo_w_PE_12_0_V_V_full_n_pass_0_in),
    .w_IO_L2_in147_U0_fifo_w_local_out_V_V_write_pass_0(w_IO_L2_in147_U0_fifo_w_local_out_V_V_write_pass_0_out),
    .cout_drain_IO_L1_out_wrapper437_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper437_U0_fifo_cout_drain_out_V_V_din_pass_0_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_4_9_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_4_9_V_V_full_n_pass_0_in),
    .cout_drain_IO_L1_out_wrapper437_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper437_U0_fifo_cout_drain_out_V_V_write_pass_0_out),
    .PE_wrapper297_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper297_U0_fifo_cout_drain_out_V_din_pass_0_in),
    .fifo_cout_drain_PE_12_3_V_full_n_pass_0(fifo_cout_drain_PE_12_3_V_full_n_pass_0_out),
    .PE_wrapper297_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper297_U0_fifo_cout_drain_out_V_write_pass_0_in),
    .PE_wrapper308_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper308_U0_fifo_w_out_V_V_din_pass_0_in),
    .fifo_w_PE_13_3_V_V_full_n_pass_0(fifo_w_PE_13_3_V_V_full_n_pass_0_out),
    .PE_wrapper308_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper308_U0_fifo_w_out_V_V_write_pass_0_in),
    .PE_wrapper296_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper296_U0_fifo_cin_out_V_V_din_pass_0_out),
    .fifo_cin_PE_13_2_V_V_full_n_pass_0(fifo_cin_PE_13_2_V_V_full_n_pass_0_in),
    .PE_wrapper296_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper296_U0_fifo_cin_out_V_V_write_pass_0_out),
    .PE_wrapper284_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper284_U0_fifo_w_out_V_V_din_pass_0_in),
    .fifo_w_PE_11_3_V_V_full_n_pass_0(fifo_w_PE_11_3_V_V_full_n_pass_0_out),
    .PE_wrapper284_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper284_U0_fifo_w_out_V_V_write_pass_0_in),
    .PE_wrapper296_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper296_U0_fifo_w_out_V_V_din_pass_0_out),
    .fifo_w_PE_12_3_V_V_full_n_pass_0(fifo_w_PE_12_3_V_V_full_n_pass_0_in),
    .PE_wrapper296_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper296_U0_fifo_w_out_V_V_write_pass_0_out),
    .PE_wrapper296_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper296_U0_fifo_cout_drain_out_V_din_pass_0_out),
    .fifo_cout_drain_PE_12_2_V_full_n_pass_0(fifo_cout_drain_PE_12_2_V_full_n_pass_0_in),
    .PE_wrapper296_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper296_U0_fifo_cout_drain_out_V_write_pass_0_out),
    .PE_wrapper262_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper262_U0_fifo_cin_out_V_V_din_pass_0_out),
    .fifo_cin_PE_10_4_V_V_full_n_pass_0(fifo_cin_PE_10_4_V_V_full_n_pass_0_in),
    .PE_wrapper262_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper262_U0_fifo_cin_out_V_V_write_pass_0_out),
    .PE_wrapper274_U0_fifo_cout_drain_out_V_din_pass_1(PE_wrapper274_U0_fifo_cout_drain_out_V_din_pass_1_in),
    .fifo_cout_drain_PE_10_4_V_full_n_pass_1(fifo_cout_drain_PE_10_4_V_full_n_pass_1_out),
    .PE_wrapper274_U0_fifo_cout_drain_out_V_write_pass_1(PE_wrapper274_U0_fifo_cout_drain_out_V_write_pass_1_in),
    .w_IO_L2_in148_U0_fifo_w_local_out_V_V_din_pass_0(w_IO_L2_in148_U0_fifo_w_local_out_V_V_din_pass_0_in),
    .fifo_w_PE_13_0_V_V_full_n_pass_0(fifo_w_PE_13_0_V_V_full_n_pass_0_out),
    .w_IO_L2_in148_U0_fifo_w_local_out_V_V_write_pass_0(w_IO_L2_in148_U0_fifo_w_local_out_V_V_write_pass_0_in),
    .cout_drain_IO_L1_out_boundary_wrapper399_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_boundary_wrapper399_U0_fifo_cout_drain_out_V_V_din_pass_0_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_2_15_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_2_15_V_V_full_n_pass_0_in),
    .cout_drain_IO_L1_out_boundary_wrapper399_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_boundary_wrapper399_U0_fifo_cout_drain_out_V_V_write_pass_0_out),
    .PE_wrapper284_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper284_U0_fifo_cin_out_V_V_din_pass_0_in),
    .fifo_cin_PE_12_2_V_V_full_n_pass_0(fifo_cin_PE_12_2_V_V_full_n_pass_0_out),
    .PE_wrapper284_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper284_U0_fifo_cin_out_V_V_write_pass_0_in),
    .cout_drain_IO_L1_out_wrapper434_U0_fifo_cout_drain_out_V_V_din_pass_1(cout_drain_IO_L1_out_wrapper434_U0_fifo_cout_drain_out_V_V_din_pass_1_in),
    .fifo_cout_drain_cout_drain_IO_L1_out_4_12_V_V_full_n_pass_1(fifo_cout_drain_cout_drain_IO_L1_out_4_12_V_V_full_n_pass_1_out),
    .cout_drain_IO_L1_out_wrapper434_U0_fifo_cout_drain_out_V_V_write_pass_1(cout_drain_IO_L1_out_wrapper434_U0_fifo_cout_drain_out_V_V_write_pass_1_in),
    .PE_wrapper285_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper285_U0_fifo_cin_out_V_V_din_pass_0_out),
    .fifo_cin_PE_12_3_V_V_full_n_pass_0(fifo_cin_PE_12_3_V_V_full_n_pass_0_in),
    .PE_wrapper285_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper285_U0_fifo_cin_out_V_V_write_pass_0_out),
    .PE_wrapper309_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper309_U0_fifo_cout_drain_out_V_din_pass_0_out),
    .fifo_cout_drain_PE_13_3_V_full_n_pass_0(fifo_cout_drain_PE_13_3_V_full_n_pass_0_in),
    .PE_wrapper309_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper309_U0_fifo_cout_drain_out_V_write_pass_0_out),
    .ap_clk(ap_clk),
    .ap_start_Boundary_X0Y4_To_X2Y4(ap_start_Boundary_X0Y4_To_X2Y4_in),
    .ap_rst_n_Boundary_X0Y4_To_X2Y4(ap_rst_n_Boundary_X0Y4_To_X2Y4_in),
    .ap_done_Boundary_X0Y4_To_X2Y4(ap_done_Boundary_X0Y4_To_X2Y4_out),
    .ap_start_Boundary_X0Y6_To_X2Y6(ap_start_Boundary_X0Y6_To_X2Y6_out),
    .ap_rst_n_Boundary_X0Y6_To_X2Y6(ap_rst_n_Boundary_X0Y6_To_X2Y6_out),
    .ap_done_Boundary_X0Y6_To_X2Y6(ap_done_Boundary_X0Y6_To_X2Y6_in)
  );


  (* keep_hierarchy = "yes" *) CR_X0Y6_To_CR_X1Y7_ctrl CR_X0Y6_To_CR_X1Y7_ctrl_U0 (
    .cout_drain_IO_L1_out_wrapper402_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper402_U0_fifo_cout_drain_out_V_V_din_pass_0_in),
    .cout_drain_IO_L1_out_wrapper402_U0_fifo_cout_drain_out_V_V_din_pass_1(cout_drain_IO_L1_out_wrapper402_U0_fifo_cout_drain_out_V_V_din_pass_1_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_2_12_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_2_12_V_V_full_n_pass_0_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_2_12_V_V_full_n_pass_1(fifo_cout_drain_cout_drain_IO_L1_out_2_12_V_V_full_n_pass_1_in),
    .cout_drain_IO_L1_out_wrapper402_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper402_U0_fifo_cout_drain_out_V_V_write_pass_0_in),
    .cout_drain_IO_L1_out_wrapper402_U0_fifo_cout_drain_out_V_V_write_pass_1(cout_drain_IO_L1_out_wrapper402_U0_fifo_cout_drain_out_V_V_write_pass_1_out),
    .PE_wrapper286_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper286_U0_fifo_cout_drain_out_V_din_pass_0_in),
    .PE_wrapper286_U0_fifo_cout_drain_out_V_din_pass_1(PE_wrapper286_U0_fifo_cout_drain_out_V_din_pass_1_out),
    .fifo_cout_drain_PE_11_4_V_full_n_pass_0(fifo_cout_drain_PE_11_4_V_full_n_pass_0_out),
    .fifo_cout_drain_PE_11_4_V_full_n_pass_1(fifo_cout_drain_PE_11_4_V_full_n_pass_1_in),
    .PE_wrapper286_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper286_U0_fifo_cout_drain_out_V_write_pass_0_in),
    .PE_wrapper286_U0_fifo_cout_drain_out_V_write_pass_1(PE_wrapper286_U0_fifo_cout_drain_out_V_write_pass_1_out),
    .PE_wrapper226_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper226_U0_fifo_cout_drain_out_V_din_pass_0_in),
    .PE_wrapper226_U0_fifo_cout_drain_out_V_din_pass_1(PE_wrapper226_U0_fifo_cout_drain_out_V_din_pass_1_out),
    .fifo_cout_drain_PE_6_4_V_full_n_pass_0(fifo_cout_drain_PE_6_4_V_full_n_pass_0_out),
    .fifo_cout_drain_PE_6_4_V_full_n_pass_1(fifo_cout_drain_PE_6_4_V_full_n_pass_1_in),
    .PE_wrapper226_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper226_U0_fifo_cout_drain_out_V_write_pass_0_in),
    .PE_wrapper226_U0_fifo_cout_drain_out_V_write_pass_1(PE_wrapper226_U0_fifo_cout_drain_out_V_write_pass_1_out),
    .PE_wrapper320_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper320_U0_fifo_cin_out_V_V_din_pass_0_in),
    .PE_wrapper320_U0_fifo_cin_out_V_V_din_pass_1(PE_wrapper320_U0_fifo_cin_out_V_V_din_pass_1_out),
    .fifo_cin_PE_15_2_V_V_full_n_pass_0(fifo_cin_PE_15_2_V_V_full_n_pass_0_out),
    .fifo_cin_PE_15_2_V_V_full_n_pass_1(fifo_cin_PE_15_2_V_V_full_n_pass_1_in),
    .PE_wrapper320_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper320_U0_fifo_cin_out_V_V_write_pass_0_in),
    .PE_wrapper320_U0_fifo_cin_out_V_V_write_pass_1(PE_wrapper320_U0_fifo_cin_out_V_V_write_pass_1_out),
    .PE_wrapper321_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper321_U0_fifo_cin_out_V_V_din_pass_0_in),
    .PE_wrapper321_U0_fifo_cin_out_V_V_din_pass_1(PE_wrapper321_U0_fifo_cin_out_V_V_din_pass_1_out),
    .fifo_cin_PE_15_3_V_V_full_n_pass_0(fifo_cin_PE_15_3_V_V_full_n_pass_0_out),
    .fifo_cin_PE_15_3_V_V_full_n_pass_1(fifo_cin_PE_15_3_V_V_full_n_pass_1_in),
    .PE_wrapper321_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper321_U0_fifo_cin_out_V_V_write_pass_0_in),
    .PE_wrapper321_U0_fifo_cin_out_V_V_write_pass_1(PE_wrapper321_U0_fifo_cin_out_V_V_write_pass_1_out),
    .PE_wrapper274_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper274_U0_fifo_cout_drain_out_V_din_pass_0_in),
    .PE_wrapper274_U0_fifo_cout_drain_out_V_din_pass_1(PE_wrapper274_U0_fifo_cout_drain_out_V_din_pass_1_out),
    .fifo_cout_drain_PE_10_4_V_full_n_pass_0(fifo_cout_drain_PE_10_4_V_full_n_pass_0_out),
    .fifo_cout_drain_PE_10_4_V_full_n_pass_1(fifo_cout_drain_PE_10_4_V_full_n_pass_1_in),
    .PE_wrapper274_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper274_U0_fifo_cout_drain_out_V_write_pass_0_in),
    .PE_wrapper274_U0_fifo_cout_drain_out_V_write_pass_1(PE_wrapper274_U0_fifo_cout_drain_out_V_write_pass_1_out),
    .cout_drain_IO_L1_out_wrapper434_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper434_U0_fifo_cout_drain_out_V_V_din_pass_0_in),
    .cout_drain_IO_L1_out_wrapper434_U0_fifo_cout_drain_out_V_V_din_pass_1(cout_drain_IO_L1_out_wrapper434_U0_fifo_cout_drain_out_V_V_din_pass_1_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_4_12_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_4_12_V_V_full_n_pass_0_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_4_12_V_V_full_n_pass_1(fifo_cout_drain_cout_drain_IO_L1_out_4_12_V_V_full_n_pass_1_in),
    .cout_drain_IO_L1_out_wrapper434_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper434_U0_fifo_cout_drain_out_V_V_write_pass_0_in),
    .cout_drain_IO_L1_out_wrapper434_U0_fifo_cout_drain_out_V_V_write_pass_1(cout_drain_IO_L1_out_wrapper434_U0_fifo_cout_drain_out_V_V_write_pass_1_out),
    .PE_wrapper262_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper262_U0_fifo_w_out_V_V_din_pass_0_in),
    .PE_wrapper262_U0_fifo_w_out_V_V_din_pass_1(PE_wrapper262_U0_fifo_w_out_V_V_din_pass_1_out),
    .fifo_w_PE_9_5_V_V_full_n_pass_0(fifo_w_PE_9_5_V_V_full_n_pass_0_out),
    .fifo_w_PE_9_5_V_V_full_n_pass_1(fifo_w_PE_9_5_V_V_full_n_pass_1_in),
    .PE_wrapper262_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper262_U0_fifo_w_out_V_V_write_pass_0_in),
    .PE_wrapper262_U0_fifo_w_out_V_V_write_pass_1(PE_wrapper262_U0_fifo_w_out_V_V_write_pass_1_out),
    .PE_wrapper298_U0_fifo_w_out_V_V_din_pass_1(PE_wrapper298_U0_fifo_w_out_V_V_din_pass_1_in),
    .PE_wrapper298_U0_fifo_w_out_V_V_din_pass_2(PE_wrapper298_U0_fifo_w_out_V_V_din_pass_2_out),
    .fifo_w_PE_12_5_V_V_full_n_pass_1(fifo_w_PE_12_5_V_V_full_n_pass_1_out),
    .fifo_w_PE_12_5_V_V_full_n_pass_2(fifo_w_PE_12_5_V_V_full_n_pass_2_in),
    .PE_wrapper298_U0_fifo_w_out_V_V_write_pass_1(PE_wrapper298_U0_fifo_w_out_V_V_write_pass_1_in),
    .PE_wrapper298_U0_fifo_w_out_V_V_write_pass_2(PE_wrapper298_U0_fifo_w_out_V_V_write_pass_2_out),
    .PE_wrapper322_U0_fifo_w_out_V_V_din_pass_1(PE_wrapper322_U0_fifo_w_out_V_V_din_pass_1_in),
    .PE_wrapper322_U0_fifo_w_out_V_V_din_pass_2(PE_wrapper322_U0_fifo_w_out_V_V_din_pass_2_out),
    .fifo_w_PE_14_5_V_V_full_n_pass_1(fifo_w_PE_14_5_V_V_full_n_pass_1_out),
    .fifo_w_PE_14_5_V_V_full_n_pass_2(fifo_w_PE_14_5_V_V_full_n_pass_2_in),
    .PE_wrapper322_U0_fifo_w_out_V_V_write_pass_1(PE_wrapper322_U0_fifo_w_out_V_V_write_pass_1_in),
    .PE_wrapper322_U0_fifo_w_out_V_V_write_pass_2(PE_wrapper322_U0_fifo_w_out_V_V_write_pass_2_out),
    .PE_wrapper334_U0_fifo_w_out_V_V_din_pass_1(PE_wrapper334_U0_fifo_w_out_V_V_din_pass_1_in),
    .PE_wrapper334_U0_fifo_w_out_V_V_din_pass_2(PE_wrapper334_U0_fifo_w_out_V_V_din_pass_2_out),
    .fifo_w_PE_15_5_V_V_full_n_pass_1(fifo_w_PE_15_5_V_V_full_n_pass_1_out),
    .fifo_w_PE_15_5_V_V_full_n_pass_2(fifo_w_PE_15_5_V_V_full_n_pass_2_in),
    .PE_wrapper334_U0_fifo_w_out_V_V_write_pass_1(PE_wrapper334_U0_fifo_w_out_V_V_write_pass_1_in),
    .PE_wrapper334_U0_fifo_w_out_V_V_write_pass_2(PE_wrapper334_U0_fifo_w_out_V_V_write_pass_2_out),
    .cout_drain_IO_L1_out_wrapper385_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper385_U0_fifo_cout_drain_out_V_V_din_pass_0_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_1_13_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_1_13_V_V_full_n_pass_0_in),
    .cout_drain_IO_L1_out_wrapper385_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper385_U0_fifo_cout_drain_out_V_V_write_pass_0_out),
    .PE_wrapper298_U0_fifo_cin_out_V_V_din_pass_1(PE_wrapper298_U0_fifo_cin_out_V_V_din_pass_1_in),
    .fifo_cin_PE_13_4_V_V_full_n_pass_1(fifo_cin_PE_13_4_V_V_full_n_pass_1_out),
    .PE_wrapper298_U0_fifo_cin_out_V_V_write_pass_1(PE_wrapper298_U0_fifo_cin_out_V_V_write_pass_1_in),
    .PE_wrapper250_U0_fifo_cout_drain_out_V_din_pass_1(PE_wrapper250_U0_fifo_cout_drain_out_V_din_pass_1_in),
    .fifo_cout_drain_PE_8_4_V_full_n_pass_1(fifo_cout_drain_PE_8_4_V_full_n_pass_1_out),
    .PE_wrapper250_U0_fifo_cout_drain_out_V_write_pass_1(PE_wrapper250_U0_fifo_cout_drain_out_V_write_pass_1_in),
    .PE_wrapper310_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper310_U0_fifo_w_out_V_V_din_pass_0_out),
    .fifo_w_PE_13_5_V_V_full_n_pass_0(fifo_w_PE_13_5_V_V_full_n_pass_0_in),
    .PE_wrapper310_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper310_U0_fifo_w_out_V_V_write_pass_0_out),
    .cout_drain_IO_L1_out_wrapper439_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper439_U0_fifo_cout_drain_out_V_V_din_pass_0_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_4_7_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_4_7_V_V_full_n_pass_0_in),
    .cout_drain_IO_L1_out_wrapper439_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper439_U0_fifo_cout_drain_out_V_V_write_pass_0_out),
    .PE_wrapper310_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper310_U0_fifo_cout_drain_out_V_din_pass_0_out),
    .fifo_cout_drain_PE_13_4_V_full_n_pass_0(fifo_cout_drain_PE_13_4_V_full_n_pass_0_in),
    .PE_wrapper310_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper310_U0_fifo_cout_drain_out_V_write_pass_0_out),
    .PE_wrapper295_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper295_U0_fifo_w_out_V_V_din_pass_0_out),
    .fifo_w_PE_12_2_V_V_full_n_pass_0(fifo_w_PE_12_2_V_V_full_n_pass_0_in),
    .PE_wrapper295_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper295_U0_fifo_w_out_V_V_write_pass_0_out),
    .w_IO_L2_in148_U0_fifo_w_out_V_V_din_pass_0(w_IO_L2_in148_U0_fifo_w_out_V_V_din_pass_0_out),
    .fifo_w_w_IO_L2_in_14_V_V_full_n_pass_0(fifo_w_w_IO_L2_in_14_V_V_full_n_pass_0_in),
    .w_IO_L2_in148_U0_fifo_w_out_V_V_write_pass_0(w_IO_L2_in148_U0_fifo_w_out_V_V_write_pass_0_out),
    .PE_wrapper309_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper309_U0_fifo_w_out_V_V_din_pass_0_in),
    .fifo_w_PE_13_4_V_V_full_n_pass_0(fifo_w_PE_13_4_V_V_full_n_pass_0_out),
    .PE_wrapper309_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper309_U0_fifo_w_out_V_V_write_pass_0_in),
    .cout_drain_IO_L1_out_wrapper417_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper417_U0_fifo_cout_drain_out_V_V_din_pass_0_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_3_13_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_3_13_V_V_full_n_pass_0_in),
    .cout_drain_IO_L1_out_wrapper417_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper417_U0_fifo_cout_drain_out_V_V_write_pass_0_out),
    .PE_wrapper308_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper308_U0_fifo_cout_drain_out_V_din_pass_0_out),
    .fifo_cout_drain_PE_13_2_V_full_n_pass_0(fifo_cout_drain_PE_13_2_V_full_n_pass_0_in),
    .PE_wrapper308_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper308_U0_fifo_cout_drain_out_V_write_pass_0_out),
    .w_IO_L2_in147_U0_fifo_w_out_V_V_din_pass_0(w_IO_L2_in147_U0_fifo_w_out_V_V_din_pass_0_in),
    .fifo_w_w_IO_L2_in_13_V_V_full_n_pass_0(fifo_w_w_IO_L2_in_13_V_V_full_n_pass_0_out),
    .w_IO_L2_in147_U0_fifo_w_out_V_V_write_pass_0(w_IO_L2_in147_U0_fifo_w_out_V_V_write_pass_0_in),
    .PE_wrapper282_U0_fifo_cin_out_V_V_din_pass_1(PE_wrapper282_U0_fifo_cin_out_V_V_din_pass_1_in),
    .fifo_cin_PE_12_0_V_V_full_n_pass_1(fifo_cin_PE_12_0_V_V_full_n_pass_1_out),
    .PE_wrapper282_U0_fifo_cin_out_V_V_write_pass_1(PE_wrapper282_U0_fifo_cin_out_V_V_write_pass_1_in),
    .cout_drain_IO_L1_out_wrapper416_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper416_U0_fifo_cout_drain_out_V_V_din_pass_0_in),
    .fifo_cout_drain_cout_drain_IO_L1_out_3_14_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_3_14_V_V_full_n_pass_0_out),
    .cout_drain_IO_L1_out_wrapper416_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper416_U0_fifo_cout_drain_out_V_V_write_pass_0_in),
    .PE_wrapper297_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper297_U0_fifo_cin_out_V_V_din_pass_0_out),
    .fifo_cin_PE_13_3_V_V_full_n_pass_0(fifo_cin_PE_13_3_V_V_full_n_pass_0_in),
    .PE_wrapper297_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper297_U0_fifo_cin_out_V_V_write_pass_0_out),
    .PE_wrapper306_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper306_U0_fifo_w_out_V_V_din_pass_0_in),
    .fifo_w_PE_13_1_V_V_full_n_pass_0(fifo_w_PE_13_1_V_V_full_n_pass_0_out),
    .PE_wrapper306_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper306_U0_fifo_w_out_V_V_write_pass_0_in),
    .PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0_out),
    .fifo_cin_PE_8_4_V_V_full_n_pass_0(fifo_cin_PE_8_4_V_V_full_n_pass_0_in),
    .PE_wrapper238_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper238_U0_fifo_cin_out_V_V_write_pass_0_out),
    .PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0_out),
    .fifo_w_PE_12_4_V_V_full_n_pass_0(fifo_w_PE_12_4_V_V_full_n_pass_0_in),
    .PE_wrapper297_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper297_U0_fifo_w_out_V_V_write_pass_0_out),
    .PE_wrapper294_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper294_U0_fifo_cout_drain_out_V_din_pass_0_out),
    .fifo_cout_drain_PE_12_0_V_full_n_pass_0(fifo_cout_drain_PE_12_0_V_full_n_pass_0_in),
    .PE_wrapper294_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper294_U0_fifo_cout_drain_out_V_write_pass_0_out),
    .PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0_out),
    .fifo_cin_PE_14_4_V_V_full_n_pass_0(fifo_cin_PE_14_4_V_V_full_n_pass_0_in),
    .PE_wrapper310_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper310_U0_fifo_cin_out_V_V_write_pass_0_out),
    .PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0_out),
    .fifo_cin_PE_14_1_V_V_full_n_pass_0(fifo_cin_PE_14_1_V_V_full_n_pass_0_in),
    .PE_wrapper307_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper307_U0_fifo_cin_out_V_V_write_pass_0_out),
    .PE_wrapper237_U0_fifo_w_out_V_V_din_pass_2(PE_wrapper237_U0_fifo_w_out_V_V_din_pass_2_in),
    .fifo_w_PE_7_4_V_V_full_n_pass_2(fifo_w_PE_7_4_V_V_full_n_pass_2_out),
    .PE_wrapper237_U0_fifo_w_out_V_V_write_pass_2(PE_wrapper237_U0_fifo_w_out_V_V_write_pass_2_in),
    .PE_wrapper283_U0_fifo_cin_out_V_V_din_pass_1(PE_wrapper283_U0_fifo_cin_out_V_V_din_pass_1_in),
    .fifo_cin_PE_12_1_V_V_full_n_pass_1(fifo_cin_PE_12_1_V_V_full_n_pass_1_out),
    .PE_wrapper283_U0_fifo_cin_out_V_V_write_pass_1(PE_wrapper283_U0_fifo_cin_out_V_V_write_pass_1_in),
    .PE_wrapper295_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper295_U0_fifo_cout_drain_out_V_din_pass_0_out),
    .fifo_cout_drain_PE_12_1_V_full_n_pass_0(fifo_cout_drain_PE_12_1_V_full_n_pass_0_in),
    .PE_wrapper295_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper295_U0_fifo_cout_drain_out_V_write_pass_0_out),
    .PE_wrapper294_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper294_U0_fifo_cin_out_V_V_din_pass_0_out),
    .fifo_cin_PE_13_0_V_V_full_n_pass_0(fifo_cin_PE_13_0_V_V_full_n_pass_0_in),
    .PE_wrapper294_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper294_U0_fifo_cin_out_V_V_write_pass_0_out),
    .w_IO_L2_in147_U0_fifo_w_local_out_V_V_din_pass_0(w_IO_L2_in147_U0_fifo_w_local_out_V_V_din_pass_0_in),
    .fifo_w_PE_12_0_V_V_full_n_pass_0(fifo_w_PE_12_0_V_V_full_n_pass_0_out),
    .w_IO_L2_in147_U0_fifo_w_local_out_V_V_write_pass_0(w_IO_L2_in147_U0_fifo_w_local_out_V_V_write_pass_0_in),
    .cout_drain_IO_L1_out_wrapper437_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper437_U0_fifo_cout_drain_out_V_V_din_pass_0_in),
    .fifo_cout_drain_cout_drain_IO_L1_out_4_9_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_4_9_V_V_full_n_pass_0_out),
    .cout_drain_IO_L1_out_wrapper437_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper437_U0_fifo_cout_drain_out_V_V_write_pass_0_in),
    .PE_wrapper297_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper297_U0_fifo_cout_drain_out_V_din_pass_0_out),
    .fifo_cout_drain_PE_12_3_V_full_n_pass_0(fifo_cout_drain_PE_12_3_V_full_n_pass_0_in),
    .PE_wrapper297_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper297_U0_fifo_cout_drain_out_V_write_pass_0_out),
    .PE_wrapper308_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper308_U0_fifo_cin_out_V_V_din_pass_0_out),
    .fifo_cin_PE_14_2_V_V_full_n_pass_0(fifo_cin_PE_14_2_V_V_full_n_pass_0_in),
    .PE_wrapper308_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper308_U0_fifo_cin_out_V_V_write_pass_0_out),
    .cout_drain_IO_L1_out_wrapper384_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper384_U0_fifo_cout_drain_out_V_V_din_pass_0_in),
    .fifo_cout_drain_cout_drain_IO_L1_out_1_14_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_1_14_V_V_full_n_pass_0_out),
    .cout_drain_IO_L1_out_wrapper384_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper384_U0_fifo_cout_drain_out_V_V_write_pass_0_in),
    .PE_wrapper308_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper308_U0_fifo_w_out_V_V_din_pass_0_out),
    .fifo_w_PE_13_3_V_V_full_n_pass_0(fifo_w_PE_13_3_V_V_full_n_pass_0_in),
    .PE_wrapper308_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper308_U0_fifo_w_out_V_V_write_pass_0_out),
    .PE_wrapper296_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper296_U0_fifo_cin_out_V_V_din_pass_0_in),
    .fifo_cin_PE_13_2_V_V_full_n_pass_0(fifo_cin_PE_13_2_V_V_full_n_pass_0_out),
    .PE_wrapper296_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper296_U0_fifo_cin_out_V_V_write_pass_0_in),
    .PE_wrapper296_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper296_U0_fifo_w_out_V_V_din_pass_0_in),
    .fifo_w_PE_12_3_V_V_full_n_pass_0(fifo_w_PE_12_3_V_V_full_n_pass_0_out),
    .PE_wrapper296_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper296_U0_fifo_w_out_V_V_write_pass_0_in),
    .PE_wrapper226_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper226_U0_fifo_cin_out_V_V_din_pass_0_in),
    .fifo_cin_PE_7_4_V_V_full_n_pass_0(fifo_cin_PE_7_4_V_V_full_n_pass_0_out),
    .PE_wrapper226_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper226_U0_fifo_cin_out_V_V_write_pass_0_in),
    .w_IO_L2_in148_U0_fifo_w_local_out_V_V_din_pass_0(w_IO_L2_in148_U0_fifo_w_local_out_V_V_din_pass_0_out),
    .fifo_w_PE_13_0_V_V_full_n_pass_0(fifo_w_PE_13_0_V_V_full_n_pass_0_in),
    .w_IO_L2_in148_U0_fifo_w_local_out_V_V_write_pass_0(w_IO_L2_in148_U0_fifo_w_local_out_V_V_write_pass_0_out),
    .PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0_out),
    .fifo_w_PE_7_5_V_V_full_n_pass_0(fifo_w_PE_7_5_V_V_full_n_pass_0_in),
    .PE_wrapper238_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper238_U0_fifo_w_out_V_V_write_pass_0_out),
    .PE_wrapper285_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper285_U0_fifo_cin_out_V_V_din_pass_0_in),
    .fifo_cin_PE_12_3_V_V_full_n_pass_0(fifo_cin_PE_12_3_V_V_full_n_pass_0_out),
    .PE_wrapper285_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper285_U0_fifo_cin_out_V_V_write_pass_0_in),
    .PE_wrapper309_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper309_U0_fifo_cout_drain_out_V_din_pass_0_in),
    .fifo_cout_drain_PE_13_3_V_full_n_pass_0(fifo_cout_drain_PE_13_3_V_full_n_pass_0_out),
    .PE_wrapper309_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper309_U0_fifo_cout_drain_out_V_write_pass_0_in),
    .ap_clk(ap_clk),
    .ap_start_Boundary_X0Y6_To_X2Y6(ap_start_Boundary_X0Y6_To_X2Y6_in),
    .ap_rst_n_Boundary_X0Y6_To_X2Y6(ap_rst_n_Boundary_X0Y6_To_X2Y6_in),
    .ap_done_Boundary_X0Y6_To_X2Y6(ap_done_Boundary_X0Y6_To_X2Y6_out),
    .ap_start_Boundary_X0Y8_To_X2Y8(ap_start_Boundary_X0Y8_To_X2Y8_out),
    .ap_rst_n_Boundary_X0Y8_To_X2Y8(ap_rst_n_Boundary_X0Y8_To_X2Y8_out),
    .ap_done_Boundary_X0Y8_To_X2Y8(ap_done_Boundary_X0Y8_To_X2Y8_in)
  );


  (* keep_hierarchy = "yes" *) CR_X2Y4_To_CR_X3Y5_ctrl CR_X2Y4_To_CR_X3Y5_ctrl_U0 (
    .PE_wrapper309_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper309_U0_fifo_cin_out_V_V_din_pass_0_in),
    .PE_wrapper309_U0_fifo_cin_out_V_V_din_pass_1(PE_wrapper309_U0_fifo_cin_out_V_V_din_pass_1_out),
    .fifo_cin_PE_14_3_V_V_full_n_pass_0(fifo_cin_PE_14_3_V_V_full_n_pass_0_out),
    .fifo_cin_PE_14_3_V_V_full_n_pass_1(fifo_cin_PE_14_3_V_V_full_n_pass_1_in),
    .PE_wrapper309_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper309_U0_fifo_cin_out_V_V_write_pass_0_in),
    .PE_wrapper309_U0_fifo_cin_out_V_V_write_pass_1(PE_wrapper309_U0_fifo_cin_out_V_V_write_pass_1_out),
    .PE_wrapper214_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper214_U0_fifo_cin_out_V_V_din_pass_0_in),
    .PE_wrapper214_U0_fifo_cin_out_V_V_din_pass_1(PE_wrapper214_U0_fifo_cin_out_V_V_din_pass_1_out),
    .fifo_cin_PE_6_4_V_V_full_n_pass_0(fifo_cin_PE_6_4_V_V_full_n_pass_0_out),
    .fifo_cin_PE_6_4_V_V_full_n_pass_1(fifo_cin_PE_6_4_V_V_full_n_pass_1_in),
    .PE_wrapper214_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper214_U0_fifo_cin_out_V_V_write_pass_0_in),
    .PE_wrapper214_U0_fifo_cin_out_V_V_write_pass_1(PE_wrapper214_U0_fifo_cin_out_V_V_write_pass_1_out),
    .cout_drain_IO_L1_out_wrapper418_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper418_U0_fifo_cout_drain_out_V_V_din_pass_0_in),
    .cout_drain_IO_L1_out_wrapper418_U0_fifo_cout_drain_out_V_V_din_pass_1(cout_drain_IO_L1_out_wrapper418_U0_fifo_cout_drain_out_V_V_din_pass_1_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_3_12_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_3_12_V_V_full_n_pass_0_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_3_12_V_V_full_n_pass_1(fifo_cout_drain_cout_drain_IO_L1_out_3_12_V_V_full_n_pass_1_in),
    .cout_drain_IO_L1_out_wrapper418_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper418_U0_fifo_cout_drain_out_V_V_write_pass_0_in),
    .cout_drain_IO_L1_out_wrapper418_U0_fifo_cout_drain_out_V_V_write_pass_1(cout_drain_IO_L1_out_wrapper418_U0_fifo_cout_drain_out_V_V_write_pass_1_out),
    .PE_wrapper225_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper225_U0_fifo_w_out_V_V_din_pass_0_in),
    .PE_wrapper225_U0_fifo_w_out_V_V_din_pass_1(PE_wrapper225_U0_fifo_w_out_V_V_din_pass_1_out),
    .fifo_w_PE_6_4_V_V_full_n_pass_0(fifo_w_PE_6_4_V_V_full_n_pass_0_out),
    .fifo_w_PE_6_4_V_V_full_n_pass_1(fifo_w_PE_6_4_V_V_full_n_pass_1_in),
    .PE_wrapper225_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper225_U0_fifo_w_out_V_V_write_pass_0_in),
    .PE_wrapper225_U0_fifo_w_out_V_V_write_pass_1(PE_wrapper225_U0_fifo_w_out_V_V_write_pass_1_out),
    .PE_wrapper285_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper285_U0_fifo_w_out_V_V_din_pass_0_in),
    .PE_wrapper285_U0_fifo_w_out_V_V_din_pass_1(PE_wrapper285_U0_fifo_w_out_V_V_din_pass_1_out),
    .fifo_w_PE_11_4_V_V_full_n_pass_0(fifo_w_PE_11_4_V_V_full_n_pass_0_out),
    .fifo_w_PE_11_4_V_V_full_n_pass_1(fifo_w_PE_11_4_V_V_full_n_pass_1_in),
    .PE_wrapper285_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper285_U0_fifo_w_out_V_V_write_pass_0_in),
    .PE_wrapper285_U0_fifo_w_out_V_V_write_pass_1(PE_wrapper285_U0_fifo_w_out_V_V_write_pass_1_out),
    .PE_wrapper306_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper306_U0_fifo_cin_out_V_V_din_pass_0_in),
    .PE_wrapper306_U0_fifo_cin_out_V_V_din_pass_1(PE_wrapper306_U0_fifo_cin_out_V_V_din_pass_1_out),
    .fifo_cin_PE_14_0_V_V_full_n_pass_0(fifo_cin_PE_14_0_V_V_full_n_pass_0_out),
    .fifo_cin_PE_14_0_V_V_full_n_pass_1(fifo_cin_PE_14_0_V_V_full_n_pass_1_in),
    .PE_wrapper306_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper306_U0_fifo_cin_out_V_V_write_pass_0_in),
    .PE_wrapper306_U0_fifo_cin_out_V_V_write_pass_1(PE_wrapper306_U0_fifo_cin_out_V_V_write_pass_1_out),
    .PE_wrapper285_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper285_U0_fifo_cout_drain_out_V_din_pass_0_in),
    .PE_wrapper285_U0_fifo_cout_drain_out_V_din_pass_1(PE_wrapper285_U0_fifo_cout_drain_out_V_din_pass_1_out),
    .fifo_cout_drain_PE_11_3_V_full_n_pass_0(fifo_cout_drain_PE_11_3_V_full_n_pass_0_out),
    .fifo_cout_drain_PE_11_3_V_full_n_pass_1(fifo_cout_drain_PE_11_3_V_full_n_pass_1_in),
    .PE_wrapper285_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper285_U0_fifo_cout_drain_out_V_write_pass_0_in),
    .PE_wrapper285_U0_fifo_cout_drain_out_V_write_pass_1(PE_wrapper285_U0_fifo_cout_drain_out_V_write_pass_1_out),
    .PE_wrapper262_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper262_U0_fifo_cin_out_V_V_din_pass_0_in),
    .PE_wrapper262_U0_fifo_cin_out_V_V_din_pass_1(PE_wrapper262_U0_fifo_cin_out_V_V_din_pass_1_out),
    .fifo_cin_PE_10_4_V_V_full_n_pass_0(fifo_cin_PE_10_4_V_V_full_n_pass_0_out),
    .fifo_cin_PE_10_4_V_V_full_n_pass_1(fifo_cin_PE_10_4_V_V_full_n_pass_1_in),
    .PE_wrapper262_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper262_U0_fifo_cin_out_V_V_write_pass_0_in),
    .PE_wrapper262_U0_fifo_cin_out_V_V_write_pass_1(PE_wrapper262_U0_fifo_cin_out_V_V_write_pass_1_out),
    .PE_wrapper296_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper296_U0_fifo_cout_drain_out_V_din_pass_0_in),
    .PE_wrapper296_U0_fifo_cout_drain_out_V_din_pass_1(PE_wrapper296_U0_fifo_cout_drain_out_V_din_pass_1_out),
    .fifo_cout_drain_PE_12_2_V_full_n_pass_0(fifo_cout_drain_PE_12_2_V_full_n_pass_0_out),
    .fifo_cout_drain_PE_12_2_V_full_n_pass_1(fifo_cout_drain_PE_12_2_V_full_n_pass_1_in),
    .PE_wrapper296_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper296_U0_fifo_cout_drain_out_V_write_pass_0_in),
    .PE_wrapper296_U0_fifo_cout_drain_out_V_write_pass_1(PE_wrapper296_U0_fifo_cout_drain_out_V_write_pass_1_out),
    .cout_drain_IO_L1_out_wrapper440_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper440_U0_fifo_cout_drain_out_V_V_din_pass_0_in),
    .cout_drain_IO_L1_out_wrapper440_U0_fifo_cout_drain_out_V_V_din_pass_1(cout_drain_IO_L1_out_wrapper440_U0_fifo_cout_drain_out_V_V_din_pass_1_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_4_6_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_4_6_V_V_full_n_pass_0_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_4_6_V_V_full_n_pass_1(fifo_cout_drain_cout_drain_IO_L1_out_4_6_V_V_full_n_pass_1_in),
    .cout_drain_IO_L1_out_wrapper440_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper440_U0_fifo_cout_drain_out_V_V_write_pass_0_in),
    .cout_drain_IO_L1_out_wrapper440_U0_fifo_cout_drain_out_V_V_write_pass_1(cout_drain_IO_L1_out_wrapper440_U0_fifo_cout_drain_out_V_V_write_pass_1_out),
    .PE_wrapper320_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper320_U0_fifo_cout_drain_out_V_din_pass_0_in),
    .fifo_cout_drain_PE_14_2_V_full_n_pass_0(fifo_cout_drain_PE_14_2_V_full_n_pass_0_out),
    .PE_wrapper320_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper320_U0_fifo_cout_drain_out_V_write_pass_0_in),
    .cout_drain_IO_L1_out_wrapper433_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper433_U0_fifo_cout_drain_out_V_V_din_pass_0_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_4_13_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_4_13_V_V_full_n_pass_0_in),
    .cout_drain_IO_L1_out_wrapper433_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper433_U0_fifo_cout_drain_out_V_V_write_pass_0_out),
    .PE_wrapper333_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper333_U0_fifo_w_out_V_V_din_pass_0_in),
    .fifo_w_PE_15_4_V_V_full_n_pass_0(fifo_w_PE_15_4_V_V_full_n_pass_0_out),
    .PE_wrapper333_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper333_U0_fifo_w_out_V_V_write_pass_0_in),
    .w_IO_L2_in149_U0_fifo_w_out_V_V_din_pass_0(w_IO_L2_in149_U0_fifo_w_out_V_V_din_pass_0_in),
    .fifo_w_w_IO_L2_in_15_V_V_full_n_pass_0(fifo_w_w_IO_L2_in_15_V_V_full_n_pass_0_out),
    .w_IO_L2_in149_U0_fifo_w_out_V_V_write_pass_0(w_IO_L2_in149_U0_fifo_w_out_V_V_write_pass_0_in),
    .PE_wrapper250_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper250_U0_fifo_cin_out_V_V_din_pass_0_out),
    .fifo_cin_PE_9_4_V_V_full_n_pass_0(fifo_cin_PE_9_4_V_V_full_n_pass_0_in),
    .PE_wrapper250_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper250_U0_fifo_cin_out_V_V_write_pass_0_out),
    .PE_wrapper250_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper250_U0_fifo_cout_drain_out_V_din_pass_0_out),
    .fifo_cout_drain_PE_8_4_V_full_n_pass_0(fifo_cout_drain_PE_8_4_V_full_n_pass_0_in),
    .PE_wrapper250_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper250_U0_fifo_cout_drain_out_V_write_pass_0_out),
    .PE_wrapper298_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper298_U0_fifo_cin_out_V_V_din_pass_0_out),
    .fifo_cin_PE_13_4_V_V_full_n_pass_0(fifo_cin_PE_13_4_V_V_full_n_pass_0_in),
    .PE_wrapper298_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper298_U0_fifo_cin_out_V_V_write_pass_0_out),
    .cout_drain_IO_L1_out_wrapper432_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper432_U0_fifo_cout_drain_out_V_V_din_pass_0_in),
    .fifo_cout_drain_cout_drain_IO_L1_out_4_14_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_4_14_V_V_full_n_pass_0_out),
    .cout_drain_IO_L1_out_wrapper432_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper432_U0_fifo_cout_drain_out_V_V_write_pass_0_in),
    .PE_wrapper318_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper318_U0_fifo_w_out_V_V_din_pass_0_in),
    .fifo_w_PE_14_1_V_V_full_n_pass_0(fifo_w_PE_14_1_V_V_full_n_pass_0_out),
    .PE_wrapper318_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper318_U0_fifo_w_out_V_V_write_pass_0_in),
    .PE_wrapper306_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper306_U0_fifo_cout_drain_out_V_din_pass_0_in),
    .fifo_cout_drain_PE_13_0_V_full_n_pass_0(fifo_cout_drain_PE_13_0_V_full_n_pass_0_out),
    .PE_wrapper306_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper306_U0_fifo_cout_drain_out_V_write_pass_0_in),
    .PE_wrapper310_U0_fifo_cout_drain_out_V_din_pass_1(PE_wrapper310_U0_fifo_cout_drain_out_V_din_pass_1_in),
    .fifo_cout_drain_PE_13_4_V_full_n_pass_1(fifo_cout_drain_PE_13_4_V_full_n_pass_1_out),
    .PE_wrapper310_U0_fifo_cout_drain_out_V_write_pass_1(PE_wrapper310_U0_fifo_cout_drain_out_V_write_pass_1_in),
    .PE_wrapper286_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper286_U0_fifo_cin_out_V_V_din_pass_0_in),
    .fifo_cin_PE_12_4_V_V_full_n_pass_0(fifo_cin_PE_12_4_V_V_full_n_pass_0_out),
    .PE_wrapper286_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper286_U0_fifo_cin_out_V_V_write_pass_0_in),
    .PE_wrapper331_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper331_U0_fifo_w_out_V_V_din_pass_0_out),
    .fifo_w_PE_15_2_V_V_full_n_pass_0(fifo_w_PE_15_2_V_V_full_n_pass_0_in),
    .PE_wrapper331_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper331_U0_fifo_w_out_V_V_write_pass_0_out),
    .PE_wrapper308_U0_fifo_cout_drain_out_V_din_pass_1(PE_wrapper308_U0_fifo_cout_drain_out_V_din_pass_1_in),
    .fifo_cout_drain_PE_13_2_V_full_n_pass_1(fifo_cout_drain_PE_13_2_V_full_n_pass_1_out),
    .PE_wrapper308_U0_fifo_cout_drain_out_V_write_pass_1(PE_wrapper308_U0_fifo_cout_drain_out_V_write_pass_1_in),
    .PE_wrapper330_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper330_U0_fifo_w_out_V_V_din_pass_0_in),
    .fifo_w_PE_15_1_V_V_full_n_pass_0(fifo_w_PE_15_1_V_V_full_n_pass_0_out),
    .PE_wrapper330_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper330_U0_fifo_w_out_V_V_write_pass_0_in),
    .PE_wrapper330_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper330_U0_fifo_cin_out_V_V_din_pass_0_in),
    .fifo_cin_PE_16_0_V_V_full_n_pass_0(fifo_cin_PE_16_0_V_V_full_n_pass_0_out),
    .PE_wrapper330_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper330_U0_fifo_cin_out_V_V_write_pass_0_in),
    .cout_drain_IO_L1_out_wrapper419_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper419_U0_fifo_cout_drain_out_V_V_din_pass_0_in),
    .fifo_cout_drain_cout_drain_IO_L1_out_3_11_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_3_11_V_V_full_n_pass_0_out),
    .cout_drain_IO_L1_out_wrapper419_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper419_U0_fifo_cout_drain_out_V_V_write_pass_0_in),
    .w_IO_L2_in_boundary_U0_fifo_w_local_out_V_V_din_pass_0(w_IO_L2_in_boundary_U0_fifo_w_local_out_V_V_din_pass_0_out),
    .fifo_w_PE_15_0_V_V_full_n_pass_0(fifo_w_PE_15_0_V_V_full_n_pass_0_in),
    .w_IO_L2_in_boundary_U0_fifo_w_local_out_V_V_write_pass_0(w_IO_L2_in_boundary_U0_fifo_w_local_out_V_V_write_pass_0_out),
    .PE_wrapper333_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper333_U0_fifo_cout_drain_out_V_din_pass_0_in),
    .fifo_cout_drain_PE_15_3_V_full_n_pass_0(fifo_cout_drain_PE_15_3_V_full_n_pass_0_out),
    .PE_wrapper333_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper333_U0_fifo_cout_drain_out_V_write_pass_0_in),
    .PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_1(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_1_in),
    .fifo_cin_PE_8_4_V_V_full_n_pass_1(fifo_cin_PE_8_4_V_V_full_n_pass_1_out),
    .PE_wrapper238_U0_fifo_cin_out_V_V_write_pass_1(PE_wrapper238_U0_fifo_cin_out_V_V_write_pass_1_in),
    .PE_wrapper297_U0_fifo_w_out_V_V_din_pass_1(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_1_in),
    .fifo_w_PE_12_4_V_V_full_n_pass_1(fifo_w_PE_12_4_V_V_full_n_pass_1_out),
    .PE_wrapper297_U0_fifo_w_out_V_V_write_pass_1(PE_wrapper297_U0_fifo_w_out_V_V_write_pass_1_in),
    .PE_wrapper273_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper273_U0_fifo_w_out_V_V_din_pass_0_out),
    .fifo_w_PE_10_4_V_V_full_n_pass_0(fifo_w_PE_10_4_V_V_full_n_pass_0_in),
    .PE_wrapper273_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper273_U0_fifo_w_out_V_V_write_pass_0_out),
    .PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_1(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_1_in),
    .fifo_cin_PE_14_4_V_V_full_n_pass_1(fifo_cin_PE_14_4_V_V_full_n_pass_1_out),
    .PE_wrapper310_U0_fifo_cin_out_V_V_write_pass_1(PE_wrapper310_U0_fifo_cin_out_V_V_write_pass_1_in),
    .cout_drain_IO_L1_out_boundary_wrapper383_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_boundary_wrapper383_U0_fifo_cout_drain_out_V_V_din_pass_0_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_1_15_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_1_15_V_V_full_n_pass_0_in),
    .cout_drain_IO_L1_out_boundary_wrapper383_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_boundary_wrapper383_U0_fifo_cout_drain_out_V_V_write_pass_0_out),
    .PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_1(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_1_in),
    .fifo_cin_PE_14_1_V_V_full_n_pass_1(fifo_cin_PE_14_1_V_V_full_n_pass_1_out),
    .PE_wrapper307_U0_fifo_cin_out_V_V_write_pass_1(PE_wrapper307_U0_fifo_cin_out_V_V_write_pass_1_in),
    .PE_wrapper330_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper330_U0_fifo_cout_drain_out_V_din_pass_0_in),
    .fifo_cout_drain_PE_15_0_V_full_n_pass_0(fifo_cout_drain_PE_15_0_V_full_n_pass_0_out),
    .PE_wrapper330_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper330_U0_fifo_cout_drain_out_V_write_pass_0_in),
    .PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0_out),
    .fifo_w_PE_8_5_V_V_full_n_pass_0(fifo_w_PE_8_5_V_V_full_n_pass_0_in),
    .PE_wrapper250_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper250_U0_fifo_w_out_V_V_write_pass_0_out),
    .PE_wrapper273_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper273_U0_fifo_cin_out_V_V_din_pass_0_out),
    .fifo_cin_PE_11_3_V_V_full_n_pass_0(fifo_cin_PE_11_3_V_V_full_n_pass_0_in),
    .PE_wrapper273_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper273_U0_fifo_cin_out_V_V_write_pass_0_out),
    .cout_drain_IO_L1_out_wrapper369_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper369_U0_fifo_cout_drain_out_V_V_din_pass_0_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_0_13_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_0_13_V_V_full_n_pass_0_in),
    .cout_drain_IO_L1_out_wrapper369_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper369_U0_fifo_cout_drain_out_V_V_write_pass_0_out),
    .PE_wrapper319_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper319_U0_fifo_w_out_V_V_din_pass_0_out),
    .fifo_w_PE_14_2_V_V_full_n_pass_0(fifo_w_PE_14_2_V_V_full_n_pass_0_in),
    .PE_wrapper319_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper319_U0_fifo_w_out_V_V_write_pass_0_out),
    .PE_wrapper249_U0_fifo_w_out_V_V_din_pass_1(PE_wrapper249_U0_fifo_w_out_V_V_din_pass_1_in),
    .fifo_w_PE_8_4_V_V_full_n_pass_1(fifo_w_PE_8_4_V_V_full_n_pass_1_out),
    .PE_wrapper249_U0_fifo_w_out_V_V_write_pass_1(PE_wrapper249_U0_fifo_w_out_V_V_write_pass_1_in),
    .PE_wrapper319_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper319_U0_fifo_cout_drain_out_V_din_pass_0_out),
    .fifo_cout_drain_PE_14_1_V_full_n_pass_0(fifo_cout_drain_PE_14_1_V_full_n_pass_0_in),
    .PE_wrapper319_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper319_U0_fifo_cout_drain_out_V_write_pass_0_out),
    .PE_wrapper298_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper298_U0_fifo_w_out_V_V_din_pass_0_out),
    .fifo_w_PE_12_5_V_V_full_n_pass_0(fifo_w_PE_12_5_V_V_full_n_pass_0_in),
    .PE_wrapper298_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper298_U0_fifo_w_out_V_V_write_pass_0_out),
    .PE_wrapper334_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper334_U0_fifo_cout_drain_out_V_din_pass_0_out),
    .fifo_cout_drain_PE_15_4_V_full_n_pass_0(fifo_cout_drain_PE_15_4_V_full_n_pass_0_in),
    .PE_wrapper334_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper334_U0_fifo_cout_drain_out_V_write_pass_0_out),
    .PE_wrapper322_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper322_U0_fifo_w_out_V_V_din_pass_0_out),
    .fifo_w_PE_14_5_V_V_full_n_pass_0(fifo_w_PE_14_5_V_V_full_n_pass_0_in),
    .PE_wrapper322_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper322_U0_fifo_w_out_V_V_write_pass_0_out),
    .cout_drain_IO_L1_out_boundary_wrapper415_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_boundary_wrapper415_U0_fifo_cout_drain_out_V_V_din_pass_0_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_3_15_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_3_15_V_V_full_n_pass_0_in),
    .cout_drain_IO_L1_out_boundary_wrapper415_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_boundary_wrapper415_U0_fifo_cout_drain_out_V_V_write_pass_0_out),
    .cout_drain_IO_L1_out_wrapper420_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper420_U0_fifo_cout_drain_out_V_V_din_pass_0_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_3_10_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_3_10_V_V_full_n_pass_0_in),
    .cout_drain_IO_L1_out_wrapper420_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper420_U0_fifo_cout_drain_out_V_V_write_pass_0_out),
    .PE_wrapper318_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper318_U0_fifo_cout_drain_out_V_din_pass_0_in),
    .fifo_cout_drain_PE_14_0_V_full_n_pass_0(fifo_cout_drain_PE_14_0_V_full_n_pass_0_out),
    .PE_wrapper318_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper318_U0_fifo_cout_drain_out_V_write_pass_0_in),
    .PE_wrapper321_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper321_U0_fifo_w_out_V_V_din_pass_0_in),
    .fifo_w_PE_14_4_V_V_full_n_pass_0(fifo_w_PE_14_4_V_V_full_n_pass_0_out),
    .PE_wrapper321_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper321_U0_fifo_w_out_V_V_write_pass_0_in),
    .PE_wrapper322_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper322_U0_fifo_cout_drain_out_V_din_pass_0_out),
    .fifo_cout_drain_PE_14_4_V_full_n_pass_0(fifo_cout_drain_PE_14_4_V_full_n_pass_0_in),
    .PE_wrapper322_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper322_U0_fifo_cout_drain_out_V_write_pass_0_out),
    .PE_wrapper334_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper334_U0_fifo_w_out_V_V_din_pass_0_out),
    .fifo_w_PE_15_5_V_V_full_n_pass_0(fifo_w_PE_15_5_V_V_full_n_pass_0_in),
    .PE_wrapper334_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper334_U0_fifo_w_out_V_V_write_pass_0_out),
    .PE_wrapper272_U0_fifo_w_out_V_V_din_pass_1(PE_wrapper272_U0_fifo_w_out_V_V_din_pass_1_in),
    .fifo_w_PE_10_3_V_V_full_n_pass_1(fifo_w_PE_10_3_V_V_full_n_pass_1_out),
    .PE_wrapper272_U0_fifo_w_out_V_V_write_pass_1(PE_wrapper272_U0_fifo_w_out_V_V_write_pass_1_in),
    .PE_wrapper261_U0_fifo_cin_out_V_V_din_pass_1(PE_wrapper261_U0_fifo_cin_out_V_V_din_pass_1_in),
    .fifo_cin_PE_10_3_V_V_full_n_pass_1(fifo_cin_PE_10_3_V_V_full_n_pass_1_out),
    .PE_wrapper261_U0_fifo_cin_out_V_V_write_pass_1(PE_wrapper261_U0_fifo_cin_out_V_V_write_pass_1_in),
    .cout_drain_IO_L1_out_boundary_wrapper399_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_boundary_wrapper399_U0_fifo_cout_drain_out_V_V_din_pass_0_in),
    .fifo_cout_drain_cout_drain_IO_L1_out_2_15_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_2_15_V_V_full_n_pass_0_out),
    .cout_drain_IO_L1_out_boundary_wrapper399_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_boundary_wrapper399_U0_fifo_cout_drain_out_V_V_write_pass_0_in),
    .cout_drain_IO_L1_out_wrapper401_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper401_U0_fifo_cout_drain_out_V_V_din_pass_0_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_2_13_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_2_13_V_V_full_n_pass_0_in),
    .cout_drain_IO_L1_out_wrapper401_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper401_U0_fifo_cout_drain_out_V_V_write_pass_0_out),
    .PE_wrapper298_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper298_U0_fifo_cout_drain_out_V_din_pass_0_out),
    .fifo_cout_drain_PE_12_4_V_full_n_pass_0(fifo_cout_drain_PE_12_4_V_full_n_pass_0_in),
    .PE_wrapper298_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper298_U0_fifo_cout_drain_out_V_write_pass_0_out),
    .ap_clk(ap_clk),
    .ap_start_Boundary_X2Y4_To_X4Y4(ap_start_Boundary_X2Y4_To_X4Y4_in),
    .ap_rst_n_Boundary_X2Y4_To_X4Y4(ap_rst_n_Boundary_X2Y4_To_X4Y4_in),
    .ap_done_Boundary_X2Y4_To_X4Y4(ap_done_Boundary_X2Y4_To_X4Y4_out),
    .ap_start_Boundary_X2Y6_To_X4Y6(ap_start_Boundary_X2Y6_To_X4Y6_out),
    .ap_rst_n_Boundary_X2Y6_To_X4Y6(ap_rst_n_Boundary_X2Y6_To_X4Y6_out),
    .ap_done_Boundary_X2Y6_To_X4Y6(ap_done_Boundary_X2Y6_To_X4Y6_in)
  );


  (* keep_hierarchy = "yes" *) CR_X2Y6_To_CR_X3Y7_ctrl CR_X2Y6_To_CR_X3Y7_ctrl_U0 (
    .PE_wrapper310_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper310_U0_fifo_cout_drain_out_V_din_pass_0_in),
    .PE_wrapper310_U0_fifo_cout_drain_out_V_din_pass_1(PE_wrapper310_U0_fifo_cout_drain_out_V_din_pass_1_out),
    .fifo_cout_drain_PE_13_4_V_full_n_pass_0(fifo_cout_drain_PE_13_4_V_full_n_pass_0_out),
    .fifo_cout_drain_PE_13_4_V_full_n_pass_1(fifo_cout_drain_PE_13_4_V_full_n_pass_1_in),
    .PE_wrapper310_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper310_U0_fifo_cout_drain_out_V_write_pass_0_in),
    .PE_wrapper310_U0_fifo_cout_drain_out_V_write_pass_1(PE_wrapper310_U0_fifo_cout_drain_out_V_write_pass_1_out),
    .PE_wrapper308_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper308_U0_fifo_cout_drain_out_V_din_pass_0_in),
    .PE_wrapper308_U0_fifo_cout_drain_out_V_din_pass_1(PE_wrapper308_U0_fifo_cout_drain_out_V_din_pass_1_out),
    .fifo_cout_drain_PE_13_2_V_full_n_pass_0(fifo_cout_drain_PE_13_2_V_full_n_pass_0_out),
    .fifo_cout_drain_PE_13_2_V_full_n_pass_1(fifo_cout_drain_PE_13_2_V_full_n_pass_1_in),
    .PE_wrapper308_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper308_U0_fifo_cout_drain_out_V_write_pass_0_in),
    .PE_wrapper308_U0_fifo_cout_drain_out_V_write_pass_1(PE_wrapper308_U0_fifo_cout_drain_out_V_write_pass_1_out),
    .PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0_in),
    .PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_1(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_1_out),
    .fifo_cin_PE_8_4_V_V_full_n_pass_0(fifo_cin_PE_8_4_V_V_full_n_pass_0_out),
    .fifo_cin_PE_8_4_V_V_full_n_pass_1(fifo_cin_PE_8_4_V_V_full_n_pass_1_in),
    .PE_wrapper238_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper238_U0_fifo_cin_out_V_V_write_pass_0_in),
    .PE_wrapper238_U0_fifo_cin_out_V_V_write_pass_1(PE_wrapper238_U0_fifo_cin_out_V_V_write_pass_1_out),
    .PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0_in),
    .PE_wrapper297_U0_fifo_w_out_V_V_din_pass_1(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_1_out),
    .fifo_w_PE_12_4_V_V_full_n_pass_0(fifo_w_PE_12_4_V_V_full_n_pass_0_out),
    .fifo_w_PE_12_4_V_V_full_n_pass_1(fifo_w_PE_12_4_V_V_full_n_pass_1_in),
    .PE_wrapper297_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper297_U0_fifo_w_out_V_V_write_pass_0_in),
    .PE_wrapper297_U0_fifo_w_out_V_V_write_pass_1(PE_wrapper297_U0_fifo_w_out_V_V_write_pass_1_out),
    .PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0_in),
    .PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_1(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_1_out),
    .fifo_cin_PE_14_4_V_V_full_n_pass_0(fifo_cin_PE_14_4_V_V_full_n_pass_0_out),
    .fifo_cin_PE_14_4_V_V_full_n_pass_1(fifo_cin_PE_14_4_V_V_full_n_pass_1_in),
    .PE_wrapper310_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper310_U0_fifo_cin_out_V_V_write_pass_0_in),
    .PE_wrapper310_U0_fifo_cin_out_V_V_write_pass_1(PE_wrapper310_U0_fifo_cin_out_V_V_write_pass_1_out),
    .PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0_in),
    .PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_1(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_1_out),
    .fifo_cin_PE_14_1_V_V_full_n_pass_0(fifo_cin_PE_14_1_V_V_full_n_pass_0_out),
    .fifo_cin_PE_14_1_V_V_full_n_pass_1(fifo_cin_PE_14_1_V_V_full_n_pass_1_in),
    .PE_wrapper307_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper307_U0_fifo_cin_out_V_V_write_pass_0_in),
    .PE_wrapper307_U0_fifo_cin_out_V_V_write_pass_1(PE_wrapper307_U0_fifo_cin_out_V_V_write_pass_1_out),
    .PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0_in),
    .PE_wrapper250_U0_fifo_w_out_V_V_din_pass_1(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_1_out),
    .fifo_w_PE_8_5_V_V_full_n_pass_0(fifo_w_PE_8_5_V_V_full_n_pass_0_out),
    .fifo_w_PE_8_5_V_V_full_n_pass_1(fifo_w_PE_8_5_V_V_full_n_pass_1_in),
    .PE_wrapper250_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper250_U0_fifo_w_out_V_V_write_pass_0_in),
    .PE_wrapper250_U0_fifo_w_out_V_V_write_pass_1(PE_wrapper250_U0_fifo_w_out_V_V_write_pass_1_out),
    .PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0_in),
    .PE_wrapper238_U0_fifo_w_out_V_V_din_pass_1(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_1_out),
    .fifo_w_PE_7_5_V_V_full_n_pass_0(fifo_w_PE_7_5_V_V_full_n_pass_0_out),
    .fifo_w_PE_7_5_V_V_full_n_pass_1(fifo_w_PE_7_5_V_V_full_n_pass_1_in),
    .PE_wrapper238_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper238_U0_fifo_w_out_V_V_write_pass_0_in),
    .PE_wrapper238_U0_fifo_w_out_V_V_write_pass_1(PE_wrapper238_U0_fifo_w_out_V_V_write_pass_1_out),
    .PE_wrapper320_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper320_U0_fifo_cout_drain_out_V_din_pass_0_out),
    .fifo_cout_drain_PE_14_2_V_full_n_pass_0(fifo_cout_drain_PE_14_2_V_full_n_pass_0_in),
    .PE_wrapper320_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper320_U0_fifo_cout_drain_out_V_write_pass_0_out),
    .cout_drain_IO_L1_out_wrapper433_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper433_U0_fifo_cout_drain_out_V_V_din_pass_0_in),
    .fifo_cout_drain_cout_drain_IO_L1_out_4_13_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_4_13_V_V_full_n_pass_0_out),
    .cout_drain_IO_L1_out_wrapper433_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper433_U0_fifo_cout_drain_out_V_V_write_pass_0_in),
    .PE_wrapper309_U0_fifo_cin_out_V_V_din_pass_1(PE_wrapper309_U0_fifo_cin_out_V_V_din_pass_1_in),
    .fifo_cin_PE_14_3_V_V_full_n_pass_1(fifo_cin_PE_14_3_V_V_full_n_pass_1_out),
    .PE_wrapper309_U0_fifo_cin_out_V_V_write_pass_1(PE_wrapper309_U0_fifo_cin_out_V_V_write_pass_1_in),
    .cout_drain_IO_L1_out_wrapper402_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper402_U0_fifo_cout_drain_out_V_V_din_pass_0_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_2_12_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_2_12_V_V_full_n_pass_0_in),
    .cout_drain_IO_L1_out_wrapper402_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper402_U0_fifo_cout_drain_out_V_V_write_pass_0_out),
    .w_IO_L2_in149_U0_fifo_w_out_V_V_din_pass_0(w_IO_L2_in149_U0_fifo_w_out_V_V_din_pass_0_out),
    .fifo_w_w_IO_L2_in_15_V_V_full_n_pass_0(fifo_w_w_IO_L2_in_15_V_V_full_n_pass_0_in),
    .w_IO_L2_in149_U0_fifo_w_out_V_V_write_pass_0(w_IO_L2_in149_U0_fifo_w_out_V_V_write_pass_0_out),
    .PE_wrapper286_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper286_U0_fifo_cout_drain_out_V_din_pass_0_out),
    .fifo_cout_drain_PE_11_4_V_full_n_pass_0(fifo_cout_drain_PE_11_4_V_full_n_pass_0_in),
    .PE_wrapper286_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper286_U0_fifo_cout_drain_out_V_write_pass_0_out),
    .PE_wrapper214_U0_fifo_cin_out_V_V_din_pass_1(PE_wrapper214_U0_fifo_cin_out_V_V_din_pass_1_in),
    .fifo_cin_PE_6_4_V_V_full_n_pass_1(fifo_cin_PE_6_4_V_V_full_n_pass_1_out),
    .PE_wrapper214_U0_fifo_cin_out_V_V_write_pass_1(PE_wrapper214_U0_fifo_cin_out_V_V_write_pass_1_in),
    .cout_drain_IO_L1_out_wrapper432_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper432_U0_fifo_cout_drain_out_V_V_din_pass_0_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_4_14_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_4_14_V_V_full_n_pass_0_in),
    .cout_drain_IO_L1_out_wrapper432_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper432_U0_fifo_cout_drain_out_V_V_write_pass_0_out),
    .PE_wrapper318_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper318_U0_fifo_w_out_V_V_din_pass_0_out),
    .fifo_w_PE_14_1_V_V_full_n_pass_0(fifo_w_PE_14_1_V_V_full_n_pass_0_in),
    .PE_wrapper318_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper318_U0_fifo_w_out_V_V_write_pass_0_out),
    .PE_wrapper226_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper226_U0_fifo_cout_drain_out_V_din_pass_0_out),
    .fifo_cout_drain_PE_6_4_V_full_n_pass_0(fifo_cout_drain_PE_6_4_V_full_n_pass_0_in),
    .PE_wrapper226_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper226_U0_fifo_cout_drain_out_V_write_pass_0_out),
    .PE_wrapper286_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper286_U0_fifo_cin_out_V_V_din_pass_0_out),
    .fifo_cin_PE_12_4_V_V_full_n_pass_0(fifo_cin_PE_12_4_V_V_full_n_pass_0_in),
    .PE_wrapper286_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper286_U0_fifo_cin_out_V_V_write_pass_0_out),
    .w_IO_L2_in148_U0_fifo_w_out_V_V_din_pass_0(w_IO_L2_in148_U0_fifo_w_out_V_V_din_pass_0_in),
    .fifo_w_w_IO_L2_in_14_V_V_full_n_pass_0(fifo_w_w_IO_L2_in_14_V_V_full_n_pass_0_out),
    .w_IO_L2_in148_U0_fifo_w_out_V_V_write_pass_0(w_IO_L2_in148_U0_fifo_w_out_V_V_write_pass_0_in),
    .PE_wrapper320_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper320_U0_fifo_cin_out_V_V_din_pass_0_out),
    .fifo_cin_PE_15_2_V_V_full_n_pass_0(fifo_cin_PE_15_2_V_V_full_n_pass_0_in),
    .PE_wrapper320_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper320_U0_fifo_cin_out_V_V_write_pass_0_out),
    .cout_drain_IO_L1_out_wrapper418_U0_fifo_cout_drain_out_V_V_din_pass_1(cout_drain_IO_L1_out_wrapper418_U0_fifo_cout_drain_out_V_V_din_pass_1_in),
    .fifo_cout_drain_cout_drain_IO_L1_out_3_12_V_V_full_n_pass_1(fifo_cout_drain_cout_drain_IO_L1_out_3_12_V_V_full_n_pass_1_out),
    .cout_drain_IO_L1_out_wrapper418_U0_fifo_cout_drain_out_V_V_write_pass_1(cout_drain_IO_L1_out_wrapper418_U0_fifo_cout_drain_out_V_V_write_pass_1_in),
    .PE_wrapper225_U0_fifo_w_out_V_V_din_pass_1(PE_wrapper225_U0_fifo_w_out_V_V_din_pass_1_in),
    .fifo_w_PE_6_4_V_V_full_n_pass_1(fifo_w_PE_6_4_V_V_full_n_pass_1_out),
    .PE_wrapper225_U0_fifo_w_out_V_V_write_pass_1(PE_wrapper225_U0_fifo_w_out_V_V_write_pass_1_in),
    .cout_drain_IO_L1_out_wrapper416_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper416_U0_fifo_cout_drain_out_V_V_din_pass_0_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_3_14_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_3_14_V_V_full_n_pass_0_in),
    .cout_drain_IO_L1_out_wrapper416_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper416_U0_fifo_cout_drain_out_V_V_write_pass_0_out),
    .PE_wrapper330_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper330_U0_fifo_cin_out_V_V_din_pass_0_out),
    .fifo_cin_PE_16_0_V_V_full_n_pass_0(fifo_cin_PE_16_0_V_V_full_n_pass_0_in),
    .PE_wrapper330_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper330_U0_fifo_cin_out_V_V_write_pass_0_out),
    .PE_wrapper330_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper330_U0_fifo_w_out_V_V_din_pass_0_out),
    .fifo_w_PE_15_1_V_V_full_n_pass_0(fifo_w_PE_15_1_V_V_full_n_pass_0_in),
    .PE_wrapper330_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper330_U0_fifo_w_out_V_V_write_pass_0_out),
    .PE_wrapper285_U0_fifo_w_out_V_V_din_pass_1(PE_wrapper285_U0_fifo_w_out_V_V_din_pass_1_in),
    .fifo_w_PE_11_4_V_V_full_n_pass_1(fifo_w_PE_11_4_V_V_full_n_pass_1_out),
    .PE_wrapper285_U0_fifo_w_out_V_V_write_pass_1(PE_wrapper285_U0_fifo_w_out_V_V_write_pass_1_in),
    .cout_drain_IO_L1_out_wrapper419_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper419_U0_fifo_cout_drain_out_V_V_din_pass_0_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_3_11_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_3_11_V_V_full_n_pass_0_in),
    .cout_drain_IO_L1_out_wrapper419_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper419_U0_fifo_cout_drain_out_V_V_write_pass_0_out),
    .w_IO_L2_in_boundary_U0_fifo_w_local_out_V_V_din_pass_0(w_IO_L2_in_boundary_U0_fifo_w_local_out_V_V_din_pass_0_in),
    .fifo_w_PE_15_0_V_V_full_n_pass_0(fifo_w_PE_15_0_V_V_full_n_pass_0_out),
    .w_IO_L2_in_boundary_U0_fifo_w_local_out_V_V_write_pass_0(w_IO_L2_in_boundary_U0_fifo_w_local_out_V_V_write_pass_0_in),
    .PE_wrapper273_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper273_U0_fifo_w_out_V_V_din_pass_0_in),
    .fifo_w_PE_10_4_V_V_full_n_pass_0(fifo_w_PE_10_4_V_V_full_n_pass_0_out),
    .PE_wrapper273_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper273_U0_fifo_w_out_V_V_write_pass_0_in),
    .PE_wrapper286_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper286_U0_fifo_w_out_V_V_din_pass_0_out),
    .fifo_w_PE_11_5_V_V_full_n_pass_0(fifo_w_PE_11_5_V_V_full_n_pass_0_in),
    .PE_wrapper286_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper286_U0_fifo_w_out_V_V_write_pass_0_out),
    .cout_drain_IO_L1_out_boundary_wrapper383_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_boundary_wrapper383_U0_fifo_cout_drain_out_V_V_din_pass_0_in),
    .fifo_cout_drain_cout_drain_IO_L1_out_1_15_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_1_15_V_V_full_n_pass_0_out),
    .cout_drain_IO_L1_out_boundary_wrapper383_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_boundary_wrapper383_U0_fifo_cout_drain_out_V_V_write_pass_0_in),
    .PE_wrapper330_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper330_U0_fifo_cout_drain_out_V_din_pass_0_out),
    .fifo_cout_drain_PE_15_0_V_full_n_pass_0(fifo_cout_drain_PE_15_0_V_full_n_pass_0_in),
    .PE_wrapper330_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper330_U0_fifo_cout_drain_out_V_write_pass_0_out),
    .PE_wrapper306_U0_fifo_cin_out_V_V_din_pass_1(PE_wrapper306_U0_fifo_cin_out_V_V_din_pass_1_in),
    .fifo_cin_PE_14_0_V_V_full_n_pass_1(fifo_cin_PE_14_0_V_V_full_n_pass_1_out),
    .PE_wrapper306_U0_fifo_cin_out_V_V_write_pass_1(PE_wrapper306_U0_fifo_cin_out_V_V_write_pass_1_in),
    .PE_wrapper321_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper321_U0_fifo_cin_out_V_V_din_pass_0_out),
    .fifo_cin_PE_15_3_V_V_full_n_pass_0(fifo_cin_PE_15_3_V_V_full_n_pass_0_in),
    .PE_wrapper321_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper321_U0_fifo_cin_out_V_V_write_pass_0_out),
    .PE_wrapper285_U0_fifo_cout_drain_out_V_din_pass_1(PE_wrapper285_U0_fifo_cout_drain_out_V_din_pass_1_in),
    .fifo_cout_drain_PE_11_3_V_full_n_pass_1(fifo_cout_drain_PE_11_3_V_full_n_pass_1_out),
    .PE_wrapper285_U0_fifo_cout_drain_out_V_write_pass_1(PE_wrapper285_U0_fifo_cout_drain_out_V_write_pass_1_in),
    .PE_wrapper319_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper319_U0_fifo_w_out_V_V_din_pass_0_in),
    .fifo_w_PE_14_2_V_V_full_n_pass_0(fifo_w_PE_14_2_V_V_full_n_pass_0_out),
    .PE_wrapper319_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper319_U0_fifo_w_out_V_V_write_pass_0_in),
    .PE_wrapper226_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper226_U0_fifo_w_out_V_V_din_pass_0_out),
    .fifo_w_PE_6_5_V_V_full_n_pass_0(fifo_w_PE_6_5_V_V_full_n_pass_0_in),
    .PE_wrapper226_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper226_U0_fifo_w_out_V_V_write_pass_0_out),
    .PE_wrapper308_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper308_U0_fifo_cin_out_V_V_din_pass_0_in),
    .fifo_cin_PE_14_2_V_V_full_n_pass_0(fifo_cin_PE_14_2_V_V_full_n_pass_0_out),
    .PE_wrapper308_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper308_U0_fifo_cin_out_V_V_write_pass_0_in),
    .cout_drain_IO_L1_out_wrapper384_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper384_U0_fifo_cout_drain_out_V_V_din_pass_0_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_1_14_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_1_14_V_V_full_n_pass_0_in),
    .cout_drain_IO_L1_out_wrapper384_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper384_U0_fifo_cout_drain_out_V_V_write_pass_0_out),
    .PE_wrapper319_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper319_U0_fifo_cout_drain_out_V_din_pass_0_in),
    .fifo_cout_drain_PE_14_1_V_full_n_pass_0(fifo_cout_drain_PE_14_1_V_full_n_pass_0_out),
    .PE_wrapper319_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper319_U0_fifo_cout_drain_out_V_write_pass_0_in),
    .PE_wrapper334_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper334_U0_fifo_cout_drain_out_V_din_pass_0_in),
    .fifo_cout_drain_PE_15_4_V_full_n_pass_0(fifo_cout_drain_PE_15_4_V_full_n_pass_0_out),
    .PE_wrapper334_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper334_U0_fifo_cout_drain_out_V_write_pass_0_in),
    .cout_drain_IO_L1_out_boundary_wrapper415_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_boundary_wrapper415_U0_fifo_cout_drain_out_V_V_din_pass_0_in),
    .fifo_cout_drain_cout_drain_IO_L1_out_3_15_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_3_15_V_V_full_n_pass_0_out),
    .cout_drain_IO_L1_out_boundary_wrapper415_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_boundary_wrapper415_U0_fifo_cout_drain_out_V_V_write_pass_0_in),
    .PE_wrapper274_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper274_U0_fifo_w_out_V_V_din_pass_0_out),
    .fifo_w_PE_10_5_V_V_full_n_pass_0(fifo_w_PE_10_5_V_V_full_n_pass_0_in),
    .PE_wrapper274_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper274_U0_fifo_w_out_V_V_write_pass_0_out),
    .PE_wrapper262_U0_fifo_cin_out_V_V_din_pass_1(PE_wrapper262_U0_fifo_cin_out_V_V_din_pass_1_in),
    .fifo_cin_PE_10_4_V_V_full_n_pass_1(fifo_cin_PE_10_4_V_V_full_n_pass_1_out),
    .PE_wrapper262_U0_fifo_cin_out_V_V_write_pass_1(PE_wrapper262_U0_fifo_cin_out_V_V_write_pass_1_in),
    .PE_wrapper226_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper226_U0_fifo_cin_out_V_V_din_pass_0_out),
    .fifo_cin_PE_7_4_V_V_full_n_pass_0(fifo_cin_PE_7_4_V_V_full_n_pass_0_in),
    .PE_wrapper226_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper226_U0_fifo_cin_out_V_V_write_pass_0_out),
    .PE_wrapper318_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper318_U0_fifo_cout_drain_out_V_din_pass_0_out),
    .fifo_cout_drain_PE_14_0_V_full_n_pass_0(fifo_cout_drain_PE_14_0_V_full_n_pass_0_in),
    .PE_wrapper318_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper318_U0_fifo_cout_drain_out_V_write_pass_0_out),
    .PE_wrapper274_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper274_U0_fifo_cout_drain_out_V_din_pass_0_out),
    .fifo_cout_drain_PE_10_4_V_full_n_pass_0(fifo_cout_drain_PE_10_4_V_full_n_pass_0_in),
    .PE_wrapper274_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper274_U0_fifo_cout_drain_out_V_write_pass_0_out),
    .PE_wrapper296_U0_fifo_cout_drain_out_V_din_pass_1(PE_wrapper296_U0_fifo_cout_drain_out_V_din_pass_1_in),
    .fifo_cout_drain_PE_12_2_V_full_n_pass_1(fifo_cout_drain_PE_12_2_V_full_n_pass_1_out),
    .PE_wrapper296_U0_fifo_cout_drain_out_V_write_pass_1(PE_wrapper296_U0_fifo_cout_drain_out_V_write_pass_1_in),
    .PE_wrapper321_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper321_U0_fifo_w_out_V_V_din_pass_0_out),
    .fifo_w_PE_14_4_V_V_full_n_pass_0(fifo_w_PE_14_4_V_V_full_n_pass_0_in),
    .PE_wrapper321_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper321_U0_fifo_w_out_V_V_write_pass_0_out),
    .PE_wrapper322_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper322_U0_fifo_cout_drain_out_V_din_pass_0_in),
    .fifo_cout_drain_PE_14_4_V_full_n_pass_0(fifo_cout_drain_PE_14_4_V_full_n_pass_0_out),
    .PE_wrapper322_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper322_U0_fifo_cout_drain_out_V_write_pass_0_in),
    .cout_drain_IO_L1_out_wrapper401_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper401_U0_fifo_cout_drain_out_V_V_din_pass_0_in),
    .fifo_cout_drain_cout_drain_IO_L1_out_2_13_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_2_13_V_V_full_n_pass_0_out),
    .cout_drain_IO_L1_out_wrapper401_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper401_U0_fifo_cout_drain_out_V_V_write_pass_0_in),
    .cout_drain_IO_L1_out_wrapper434_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper434_U0_fifo_cout_drain_out_V_V_din_pass_0_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_4_12_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_4_12_V_V_full_n_pass_0_in),
    .cout_drain_IO_L1_out_wrapper434_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper434_U0_fifo_cout_drain_out_V_V_write_pass_0_out),
    .PE_wrapper298_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper298_U0_fifo_cout_drain_out_V_din_pass_0_in),
    .fifo_cout_drain_PE_12_4_V_full_n_pass_0(fifo_cout_drain_PE_12_4_V_full_n_pass_0_out),
    .PE_wrapper298_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper298_U0_fifo_cout_drain_out_V_write_pass_0_in),
    .ap_clk(ap_clk),
    .ap_start_Boundary_X2Y6_To_X4Y6(ap_start_Boundary_X2Y6_To_X4Y6_in),
    .ap_rst_n_Boundary_X2Y6_To_X4Y6(ap_rst_n_Boundary_X2Y6_To_X4Y6_in),
    .ap_done_Boundary_X2Y6_To_X4Y6(ap_done_Boundary_X2Y6_To_X4Y6_out),
    .ap_start_Boundary_X2Y8_To_X4Y8(ap_start_Boundary_X2Y8_To_X4Y8_out),
    .ap_rst_n_Boundary_X2Y8_To_X4Y8(ap_rst_n_Boundary_X2Y8_To_X4Y8_out),
    .ap_done_Boundary_X2Y8_To_X4Y8(ap_done_Boundary_X2Y8_To_X4Y8_in)
  );


  (* keep_hierarchy = "yes" *) CR_X0Y8_To_CR_X1Y9_ctrl CR_X0Y8_To_CR_X1Y9_ctrl_U0 (
    .PE_wrapper288_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper288_U0_fifo_cin_out_V_V_din_pass_0_in),
    .PE_wrapper288_U0_fifo_cin_out_V_V_din_pass_1(PE_wrapper288_U0_fifo_cin_out_V_V_din_pass_1_out),
    .fifo_cin_PE_12_6_V_V_full_n_pass_0(fifo_cin_PE_12_6_V_V_full_n_pass_0_out),
    .fifo_cin_PE_12_6_V_V_full_n_pass_1(fifo_cin_PE_12_6_V_V_full_n_pass_1_in),
    .PE_wrapper288_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper288_U0_fifo_cin_out_V_V_write_pass_0_in),
    .PE_wrapper288_U0_fifo_cin_out_V_V_write_pass_1(PE_wrapper288_U0_fifo_cin_out_V_V_write_pass_1_out),
    .PE_wrapper311_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper311_U0_fifo_w_out_V_V_din_pass_0_out),
    .fifo_w_PE_13_6_V_V_full_n_pass_0(fifo_w_PE_13_6_V_V_full_n_pass_0_in),
    .PE_wrapper311_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper311_U0_fifo_w_out_V_V_write_pass_0_out),
    .PE_wrapper251_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper251_U0_fifo_cin_out_V_V_din_pass_0_in),
    .fifo_cin_PE_9_5_V_V_full_n_pass_0(fifo_cin_PE_9_5_V_V_full_n_pass_0_out),
    .PE_wrapper251_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper251_U0_fifo_cin_out_V_V_write_pass_0_in),
    .PE_wrapper299_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper299_U0_fifo_w_out_V_V_din_pass_0_out),
    .fifo_w_PE_12_6_V_V_full_n_pass_0(fifo_w_PE_12_6_V_V_full_n_pass_0_in),
    .PE_wrapper299_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper299_U0_fifo_w_out_V_V_write_pass_0_out),
    .PE_wrapper263_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper263_U0_fifo_cout_drain_out_V_din_pass_0_out),
    .fifo_cout_drain_PE_9_5_V_full_n_pass_0(fifo_cout_drain_PE_9_5_V_full_n_pass_0_in),
    .PE_wrapper263_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper263_U0_fifo_cout_drain_out_V_write_pass_0_out),
    .PE_wrapper310_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper310_U0_fifo_w_out_V_V_din_pass_0_in),
    .fifo_w_PE_13_5_V_V_full_n_pass_0(fifo_w_PE_13_5_V_V_full_n_pass_0_out),
    .PE_wrapper310_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper310_U0_fifo_w_out_V_V_write_pass_0_in),
    .PE_wrapper336_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper336_U0_fifo_cout_drain_out_V_din_pass_0_out),
    .fifo_cout_drain_PE_15_6_V_full_n_pass_0(fifo_cout_drain_PE_15_6_V_full_n_pass_0_in),
    .PE_wrapper336_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper336_U0_fifo_cout_drain_out_V_write_pass_0_out),
    .PE_wrapper262_U0_fifo_w_out_V_V_din_pass_1(PE_wrapper262_U0_fifo_w_out_V_V_din_pass_1_in),
    .fifo_w_PE_9_5_V_V_full_n_pass_1(fifo_w_PE_9_5_V_V_full_n_pass_1_out),
    .PE_wrapper262_U0_fifo_w_out_V_V_write_pass_1(PE_wrapper262_U0_fifo_w_out_V_V_write_pass_1_in),
    .PE_wrapper337_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper337_U0_fifo_w_out_V_V_din_pass_0_out),
    .fifo_w_PE_15_8_V_V_full_n_pass_0(fifo_w_PE_15_8_V_V_full_n_pass_0_in),
    .PE_wrapper337_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper337_U0_fifo_w_out_V_V_write_pass_0_out),
    .cout_drain_IO_L1_out_wrapper450_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper450_U0_fifo_cout_drain_out_V_V_din_pass_0_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_5_12_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_5_12_V_V_full_n_pass_0_in),
    .cout_drain_IO_L1_out_wrapper450_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper450_U0_fifo_cout_drain_out_V_V_write_pass_0_out),
    .PE_wrapper298_U0_fifo_w_out_V_V_din_pass_2(PE_wrapper298_U0_fifo_w_out_V_V_din_pass_2_in),
    .fifo_w_PE_12_5_V_V_full_n_pass_2(fifo_w_PE_12_5_V_V_full_n_pass_2_out),
    .PE_wrapper298_U0_fifo_w_out_V_V_write_pass_2(PE_wrapper298_U0_fifo_w_out_V_V_write_pass_2_in),
    .PE_wrapper322_U0_fifo_w_out_V_V_din_pass_2(PE_wrapper322_U0_fifo_w_out_V_V_din_pass_2_in),
    .fifo_w_PE_14_5_V_V_full_n_pass_2(fifo_w_PE_14_5_V_V_full_n_pass_2_out),
    .PE_wrapper322_U0_fifo_w_out_V_V_write_pass_2(PE_wrapper322_U0_fifo_w_out_V_V_write_pass_2_in),
    .PE_wrapper263_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper263_U0_fifo_w_out_V_V_din_pass_0_out),
    .fifo_w_PE_9_6_V_V_full_n_pass_0(fifo_w_PE_9_6_V_V_full_n_pass_0_in),
    .PE_wrapper263_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper263_U0_fifo_w_out_V_V_write_pass_0_out),
    .PE_wrapper323_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper323_U0_fifo_w_out_V_V_din_pass_0_out),
    .fifo_w_PE_14_6_V_V_full_n_pass_0(fifo_w_PE_14_6_V_V_full_n_pass_0_in),
    .PE_wrapper323_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper323_U0_fifo_w_out_V_V_write_pass_0_out),
    .PE_wrapper337_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper337_U0_fifo_cout_drain_out_V_din_pass_0_out),
    .fifo_cout_drain_PE_15_7_V_full_n_pass_0(fifo_cout_drain_PE_15_7_V_full_n_pass_0_in),
    .PE_wrapper337_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper337_U0_fifo_cout_drain_out_V_write_pass_0_out),
    .PE_wrapper324_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper324_U0_fifo_cin_out_V_V_din_pass_0_in),
    .fifo_cin_PE_15_6_V_V_full_n_pass_0(fifo_cin_PE_15_6_V_V_full_n_pass_0_out),
    .PE_wrapper324_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper324_U0_fifo_cin_out_V_V_write_pass_0_in),
    .PE_wrapper334_U0_fifo_w_out_V_V_din_pass_2(PE_wrapper334_U0_fifo_w_out_V_V_din_pass_2_in),
    .fifo_w_PE_15_5_V_V_full_n_pass_2(fifo_w_PE_15_5_V_V_full_n_pass_2_out),
    .PE_wrapper334_U0_fifo_w_out_V_V_write_pass_2(PE_wrapper334_U0_fifo_w_out_V_V_write_pass_2_in),
    .PE_wrapper263_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper263_U0_fifo_cin_out_V_V_din_pass_0_out),
    .fifo_cin_PE_10_5_V_V_full_n_pass_0(fifo_cin_PE_10_5_V_V_full_n_pass_0_in),
    .PE_wrapper263_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper263_U0_fifo_cin_out_V_V_write_pass_0_out),
    .PE_wrapper325_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper325_U0_fifo_cin_out_V_V_din_pass_0_in),
    .fifo_cin_PE_15_7_V_V_full_n_pass_0(fifo_cin_PE_15_7_V_V_full_n_pass_0_out),
    .PE_wrapper325_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper325_U0_fifo_cin_out_V_V_write_pass_0_in),
    .PE_wrapper287_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper287_U0_fifo_cin_out_V_V_din_pass_0_in),
    .fifo_cin_PE_12_5_V_V_full_n_pass_0(fifo_cin_PE_12_5_V_V_full_n_pass_0_out),
    .PE_wrapper287_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper287_U0_fifo_cin_out_V_V_write_pass_0_in),
    .ap_clk(ap_clk),
    .ap_start_Boundary_X0Y8_To_X2Y8(ap_start_Boundary_X0Y8_To_X2Y8_in),
    .ap_rst_n_Boundary_X0Y8_To_X2Y8(ap_rst_n_Boundary_X0Y8_To_X2Y8_in),
    .ap_done_Boundary_X0Y8_To_X2Y8(ap_done_Boundary_X0Y8_To_X2Y8_out),
    .ap_start_Boundary_X0Y10_To_X2Y10(ap_start_Boundary_X0Y10_To_X2Y10_out),
    .ap_rst_n_Boundary_X0Y10_To_X2Y10(ap_rst_n_Boundary_X0Y10_To_X2Y10_out),
    .ap_done_Boundary_X0Y10_To_X2Y10(ap_done_Boundary_X0Y10_To_X2Y10_in)
  );


  (* keep_hierarchy = "yes" *) CR_X0Y10_To_CR_X1Y11_ctrl CR_X0Y10_To_CR_X1Y11_ctrl_U0 (
    .PE_wrapper337_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper337_U0_fifo_w_out_V_V_din_pass_0_in),
    .PE_wrapper337_U0_fifo_w_out_V_V_din_pass_1(PE_wrapper337_U0_fifo_w_out_V_V_din_pass_1_out),
    .fifo_w_PE_15_8_V_V_full_n_pass_0(fifo_w_PE_15_8_V_V_full_n_pass_0_out),
    .fifo_w_PE_15_8_V_V_full_n_pass_1(fifo_w_PE_15_8_V_V_full_n_pass_1_in),
    .PE_wrapper337_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper337_U0_fifo_w_out_V_V_write_pass_0_in),
    .PE_wrapper337_U0_fifo_w_out_V_V_write_pass_1(PE_wrapper337_U0_fifo_w_out_V_V_write_pass_1_out),
    .PE_wrapper311_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper311_U0_fifo_w_out_V_V_din_pass_0_in),
    .fifo_w_PE_13_6_V_V_full_n_pass_0(fifo_w_PE_13_6_V_V_full_n_pass_0_out),
    .PE_wrapper311_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper311_U0_fifo_w_out_V_V_write_pass_0_in),
    .PE_wrapper299_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper299_U0_fifo_w_out_V_V_din_pass_0_in),
    .fifo_w_PE_12_6_V_V_full_n_pass_0(fifo_w_PE_12_6_V_V_full_n_pass_0_out),
    .PE_wrapper299_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper299_U0_fifo_w_out_V_V_write_pass_0_in),
    .PE_wrapper289_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper289_U0_fifo_cin_out_V_V_din_pass_0_in),
    .fifo_cin_PE_12_7_V_V_full_n_pass_0(fifo_cin_PE_12_7_V_V_full_n_pass_0_out),
    .PE_wrapper289_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper289_U0_fifo_cin_out_V_V_write_pass_0_in),
    .cout_drain_IO_L1_out_wrapper466_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper466_U0_fifo_cout_drain_out_V_V_din_pass_0_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_6_12_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_6_12_V_V_full_n_pass_0_in),
    .cout_drain_IO_L1_out_wrapper466_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper466_U0_fifo_cout_drain_out_V_V_write_pass_0_out),
    .PE_wrapper290_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper290_U0_fifo_cin_out_V_V_din_pass_0_in),
    .fifo_cin_PE_12_8_V_V_full_n_pass_0(fifo_cin_PE_12_8_V_V_full_n_pass_0_out),
    .PE_wrapper290_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper290_U0_fifo_cin_out_V_V_write_pass_0_in),
    .PE_wrapper302_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper302_U0_fifo_w_out_V_V_din_pass_0_out),
    .fifo_w_PE_12_9_V_V_full_n_pass_0(fifo_w_PE_12_9_V_V_full_n_pass_0_in),
    .PE_wrapper302_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper302_U0_fifo_w_out_V_V_write_pass_0_out),
    .PE_wrapper325_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper325_U0_fifo_w_out_V_V_din_pass_0_out),
    .fifo_w_PE_14_8_V_V_full_n_pass_0(fifo_w_PE_14_8_V_V_full_n_pass_0_in),
    .PE_wrapper325_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper325_U0_fifo_w_out_V_V_write_pass_0_out),
    .PE_wrapper336_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper336_U0_fifo_cout_drain_out_V_din_pass_0_in),
    .fifo_cout_drain_PE_15_6_V_full_n_pass_0(fifo_cout_drain_PE_15_6_V_full_n_pass_0_out),
    .PE_wrapper336_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper336_U0_fifo_cout_drain_out_V_write_pass_0_in),
    .PE_wrapper302_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper302_U0_fifo_cout_drain_out_V_din_pass_0_out),
    .fifo_cout_drain_PE_12_8_V_full_n_pass_0(fifo_cout_drain_PE_12_8_V_full_n_pass_0_in),
    .PE_wrapper302_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper302_U0_fifo_cout_drain_out_V_write_pass_0_out),
    .PE_wrapper302_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper302_U0_fifo_cin_out_V_V_din_pass_0_out),
    .fifo_cin_PE_13_8_V_V_full_n_pass_0(fifo_cin_PE_13_8_V_V_full_n_pass_0_in),
    .PE_wrapper302_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper302_U0_fifo_cin_out_V_V_write_pass_0_out),
    .PE_wrapper288_U0_fifo_cin_out_V_V_din_pass_1(PE_wrapper288_U0_fifo_cin_out_V_V_din_pass_1_in),
    .fifo_cin_PE_12_6_V_V_full_n_pass_1(fifo_cin_PE_12_6_V_V_full_n_pass_1_out),
    .PE_wrapper288_U0_fifo_cin_out_V_V_write_pass_1(PE_wrapper288_U0_fifo_cin_out_V_V_write_pass_1_in),
    .PE_wrapper323_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper323_U0_fifo_w_out_V_V_din_pass_0_in),
    .fifo_w_PE_14_6_V_V_full_n_pass_0(fifo_w_PE_14_6_V_V_full_n_pass_0_out),
    .PE_wrapper323_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper323_U0_fifo_w_out_V_V_write_pass_0_in),
    .PE_wrapper337_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper337_U0_fifo_cout_drain_out_V_din_pass_0_in),
    .fifo_cout_drain_PE_15_7_V_full_n_pass_0(fifo_cout_drain_PE_15_7_V_full_n_pass_0_out),
    .PE_wrapper337_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper337_U0_fifo_cout_drain_out_V_write_pass_0_in),
    .PE_wrapper324_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper324_U0_fifo_cin_out_V_V_din_pass_0_out),
    .fifo_cin_PE_15_6_V_V_full_n_pass_0(fifo_cin_PE_15_6_V_V_full_n_pass_0_in),
    .PE_wrapper324_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper324_U0_fifo_cin_out_V_V_write_pass_0_out),
    .PE_wrapper313_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper313_U0_fifo_w_out_V_V_din_pass_0_out),
    .fifo_w_PE_13_8_V_V_full_n_pass_0(fifo_w_PE_13_8_V_V_full_n_pass_0_in),
    .PE_wrapper313_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper313_U0_fifo_w_out_V_V_write_pass_0_out),
    .PE_wrapper325_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper325_U0_fifo_cin_out_V_V_din_pass_0_out),
    .fifo_cin_PE_15_7_V_V_full_n_pass_0(fifo_cin_PE_15_7_V_V_full_n_pass_0_in),
    .PE_wrapper325_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper325_U0_fifo_cin_out_V_V_write_pass_0_out),
    .cout_drain_IO_L1_out_wrapper482_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper482_U0_fifo_cout_drain_out_V_V_din_pass_0_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_7_12_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_7_12_V_V_full_n_pass_0_in),
    .cout_drain_IO_L1_out_wrapper482_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper482_U0_fifo_cout_drain_out_V_V_write_pass_0_out),
    .ap_clk(ap_clk),
    .ap_start_Boundary_X0Y10_To_X2Y10(ap_start_Boundary_X0Y10_To_X2Y10_in),
    .ap_rst_n_Boundary_X0Y10_To_X2Y10(ap_rst_n_Boundary_X0Y10_To_X2Y10_in),
    .ap_done_Boundary_X0Y10_To_X2Y10(ap_done_Boundary_X0Y10_To_X2Y10_out),
    .ap_start_Boundary_X0Y12_To_X2Y12(ap_start_Boundary_X0Y12_To_X2Y12_out),
    .ap_rst_n_Boundary_X0Y12_To_X2Y12(ap_rst_n_Boundary_X0Y12_To_X2Y12_out),
    .ap_done_Boundary_X0Y12_To_X2Y12(ap_done_Boundary_X0Y12_To_X2Y12_in)
  );


  (* keep_hierarchy = "yes" *) CR_X2Y8_To_CR_X3Y9_ctrl CR_X2Y8_To_CR_X3Y9_ctrl_U0 (
    .PE_wrapper263_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper263_U0_fifo_w_out_V_V_din_pass_0_in),
    .PE_wrapper263_U0_fifo_w_out_V_V_din_pass_1(PE_wrapper263_U0_fifo_w_out_V_V_din_pass_1_out),
    .fifo_w_PE_9_6_V_V_full_n_pass_0(fifo_w_PE_9_6_V_V_full_n_pass_0_out),
    .fifo_w_PE_9_6_V_V_full_n_pass_1(fifo_w_PE_9_6_V_V_full_n_pass_1_in),
    .PE_wrapper263_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper263_U0_fifo_w_out_V_V_write_pass_0_in),
    .PE_wrapper263_U0_fifo_w_out_V_V_write_pass_1(PE_wrapper263_U0_fifo_w_out_V_V_write_pass_1_out),
    .PE_wrapper251_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper251_U0_fifo_cin_out_V_V_din_pass_0_out),
    .fifo_cin_PE_9_5_V_V_full_n_pass_0(fifo_cin_PE_9_5_V_V_full_n_pass_0_in),
    .PE_wrapper251_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper251_U0_fifo_cin_out_V_V_write_pass_0_out),
    .PE_wrapper263_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper263_U0_fifo_cout_drain_out_V_din_pass_0_in),
    .fifo_cout_drain_PE_9_5_V_full_n_pass_0(fifo_cout_drain_PE_9_5_V_full_n_pass_0_out),
    .PE_wrapper263_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper263_U0_fifo_cout_drain_out_V_write_pass_0_in),
    .PE_wrapper276_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper276_U0_fifo_w_out_V_V_din_pass_0_out),
    .fifo_w_PE_10_7_V_V_full_n_pass_0(fifo_w_PE_10_7_V_V_full_n_pass_0_in),
    .PE_wrapper276_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper276_U0_fifo_w_out_V_V_write_pass_0_out),
    .PE_wrapper264_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper264_U0_fifo_cout_drain_out_V_din_pass_0_in),
    .fifo_cout_drain_PE_9_6_V_full_n_pass_0(fifo_cout_drain_PE_9_6_V_full_n_pass_0_out),
    .PE_wrapper264_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper264_U0_fifo_cout_drain_out_V_write_pass_0_in),
    .cout_drain_IO_L1_out_wrapper466_U0_fifo_cout_drain_out_V_V_din_pass_1(cout_drain_IO_L1_out_wrapper466_U0_fifo_cout_drain_out_V_V_din_pass_1_in),
    .fifo_cout_drain_cout_drain_IO_L1_out_6_12_V_V_full_n_pass_1(fifo_cout_drain_cout_drain_IO_L1_out_6_12_V_V_full_n_pass_1_out),
    .cout_drain_IO_L1_out_wrapper466_U0_fifo_cout_drain_out_V_V_write_pass_1(cout_drain_IO_L1_out_wrapper466_U0_fifo_cout_drain_out_V_V_write_pass_1_in),
    .PE_wrapper264_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper264_U0_fifo_cin_out_V_V_din_pass_0_in),
    .fifo_cin_PE_10_6_V_V_full_n_pass_0(fifo_cin_PE_10_6_V_V_full_n_pass_0_out),
    .PE_wrapper264_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper264_U0_fifo_cin_out_V_V_write_pass_0_in),
    .PE_wrapper286_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper286_U0_fifo_w_out_V_V_din_pass_0_in),
    .fifo_w_PE_11_5_V_V_full_n_pass_0(fifo_w_PE_11_5_V_V_full_n_pass_0_out),
    .PE_wrapper286_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper286_U0_fifo_w_out_V_V_write_pass_0_in),
    .PE_wrapper215_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper215_U0_fifo_cin_out_V_V_din_pass_0_in),
    .fifo_cin_PE_6_5_V_V_full_n_pass_0(fifo_cin_PE_6_5_V_V_full_n_pass_0_out),
    .PE_wrapper215_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper215_U0_fifo_cin_out_V_V_write_pass_0_in),
    .PE_wrapper227_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper227_U0_fifo_w_out_V_V_din_pass_0_out),
    .fifo_w_PE_6_6_V_V_full_n_pass_0(fifo_w_PE_6_6_V_V_full_n_pass_0_in),
    .PE_wrapper227_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper227_U0_fifo_w_out_V_V_write_pass_0_out),
    .PE_wrapper250_U0_fifo_w_out_V_V_din_pass_1(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_1_in),
    .fifo_w_PE_8_5_V_V_full_n_pass_1(fifo_w_PE_8_5_V_V_full_n_pass_1_out),
    .PE_wrapper250_U0_fifo_w_out_V_V_write_pass_1(PE_wrapper250_U0_fifo_w_out_V_V_write_pass_1_in),
    .cout_drain_IO_L1_out_wrapper450_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper450_U0_fifo_cout_drain_out_V_V_din_pass_0_in),
    .fifo_cout_drain_cout_drain_IO_L1_out_5_12_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_5_12_V_V_full_n_pass_0_out),
    .cout_drain_IO_L1_out_wrapper450_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper450_U0_fifo_cout_drain_out_V_V_write_pass_0_in),
    .PE_wrapper226_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper226_U0_fifo_w_out_V_V_din_pass_0_in),
    .fifo_w_PE_6_5_V_V_full_n_pass_0(fifo_w_PE_6_5_V_V_full_n_pass_0_out),
    .PE_wrapper226_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper226_U0_fifo_w_out_V_V_write_pass_0_in),
    .cout_drain_IO_L1_out_wrapper456_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper456_U0_fifo_cout_drain_out_V_V_din_pass_0_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_5_6_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_5_6_V_V_full_n_pass_0_in),
    .cout_drain_IO_L1_out_wrapper456_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper456_U0_fifo_cout_drain_out_V_V_write_pass_0_out),
    .PE_wrapper288_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper288_U0_fifo_cin_out_V_V_din_pass_0_out),
    .fifo_cin_PE_12_6_V_V_full_n_pass_0(fifo_cin_PE_12_6_V_V_full_n_pass_0_in),
    .PE_wrapper288_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper288_U0_fifo_cin_out_V_V_write_pass_0_out),
    .PE_wrapper251_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper251_U0_fifo_w_out_V_V_din_pass_0_out),
    .fifo_w_PE_8_6_V_V_full_n_pass_0(fifo_w_PE_8_6_V_V_full_n_pass_0_in),
    .PE_wrapper251_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper251_U0_fifo_w_out_V_V_write_pass_0_out),
    .PE_wrapper274_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper274_U0_fifo_w_out_V_V_din_pass_0_in),
    .fifo_w_PE_10_5_V_V_full_n_pass_0(fifo_w_PE_10_5_V_V_full_n_pass_0_out),
    .PE_wrapper274_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper274_U0_fifo_w_out_V_V_write_pass_0_in),
    .PE_wrapper239_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper239_U0_fifo_w_out_V_V_din_pass_0_out),
    .fifo_w_PE_7_6_V_V_full_n_pass_0(fifo_w_PE_7_6_V_V_full_n_pass_0_in),
    .PE_wrapper239_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper239_U0_fifo_w_out_V_V_write_pass_0_out),
    .PE_wrapper238_U0_fifo_w_out_V_V_din_pass_1(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_1_in),
    .fifo_w_PE_7_5_V_V_full_n_pass_1(fifo_w_PE_7_5_V_V_full_n_pass_1_out),
    .PE_wrapper238_U0_fifo_w_out_V_V_write_pass_1(PE_wrapper238_U0_fifo_w_out_V_V_write_pass_1_in),
    .PE_wrapper263_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper263_U0_fifo_cin_out_V_V_din_pass_0_in),
    .fifo_cin_PE_10_5_V_V_full_n_pass_0(fifo_cin_PE_10_5_V_V_full_n_pass_0_out),
    .PE_wrapper263_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper263_U0_fifo_cin_out_V_V_write_pass_0_in),
    .cout_drain_IO_L1_out_wrapper469_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper469_U0_fifo_cout_drain_out_V_V_din_pass_0_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_6_9_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_6_9_V_V_full_n_pass_0_in),
    .cout_drain_IO_L1_out_wrapper469_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper469_U0_fifo_cout_drain_out_V_V_write_pass_0_out),
    .PE_wrapper288_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper288_U0_fifo_w_out_V_V_din_pass_0_out),
    .fifo_w_PE_11_7_V_V_full_n_pass_0(fifo_w_PE_11_7_V_V_full_n_pass_0_in),
    .PE_wrapper288_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper288_U0_fifo_w_out_V_V_write_pass_0_out),
    .PE_wrapper287_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper287_U0_fifo_cin_out_V_V_din_pass_0_out),
    .fifo_cin_PE_12_5_V_V_full_n_pass_0(fifo_cin_PE_12_5_V_V_full_n_pass_0_in),
    .PE_wrapper287_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper287_U0_fifo_cin_out_V_V_write_pass_0_out),
    .ap_clk(ap_clk),
    .ap_start_Boundary_X2Y8_To_X4Y8(ap_start_Boundary_X2Y8_To_X4Y8_in),
    .ap_rst_n_Boundary_X2Y8_To_X4Y8(ap_rst_n_Boundary_X2Y8_To_X4Y8_in),
    .ap_done_Boundary_X2Y8_To_X4Y8(ap_done_Boundary_X2Y8_To_X4Y8_out),
    .ap_start_Boundary_X2Y10_To_X4Y10(ap_start_Boundary_X2Y10_To_X4Y10_out),
    .ap_rst_n_Boundary_X2Y10_To_X4Y10(ap_rst_n_Boundary_X2Y10_To_X4Y10_out),
    .ap_done_Boundary_X2Y10_To_X4Y10(ap_done_Boundary_X2Y10_To_X4Y10_in)
  );


  (* keep_hierarchy = "yes" *) CR_X2Y10_To_CR_X3Y11_ctrl CR_X2Y10_To_CR_X3Y11_ctrl_U0 (
    .cout_drain_IO_L1_out_wrapper466_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper466_U0_fifo_cout_drain_out_V_V_din_pass_0_in),
    .cout_drain_IO_L1_out_wrapper466_U0_fifo_cout_drain_out_V_V_din_pass_1(cout_drain_IO_L1_out_wrapper466_U0_fifo_cout_drain_out_V_V_din_pass_1_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_6_12_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_6_12_V_V_full_n_pass_0_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_6_12_V_V_full_n_pass_1(fifo_cout_drain_cout_drain_IO_L1_out_6_12_V_V_full_n_pass_1_in),
    .cout_drain_IO_L1_out_wrapper466_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper466_U0_fifo_cout_drain_out_V_V_write_pass_0_in),
    .cout_drain_IO_L1_out_wrapper466_U0_fifo_cout_drain_out_V_V_write_pass_1(cout_drain_IO_L1_out_wrapper466_U0_fifo_cout_drain_out_V_V_write_pass_1_out),
    .PE_wrapper302_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper302_U0_fifo_w_out_V_V_din_pass_0_in),
    .PE_wrapper302_U0_fifo_w_out_V_V_din_pass_1(PE_wrapper302_U0_fifo_w_out_V_V_din_pass_1_out),
    .fifo_w_PE_12_9_V_V_full_n_pass_0(fifo_w_PE_12_9_V_V_full_n_pass_0_out),
    .fifo_w_PE_12_9_V_V_full_n_pass_1(fifo_w_PE_12_9_V_V_full_n_pass_1_in),
    .PE_wrapper302_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper302_U0_fifo_w_out_V_V_write_pass_0_in),
    .PE_wrapper302_U0_fifo_w_out_V_V_write_pass_1(PE_wrapper302_U0_fifo_w_out_V_V_write_pass_1_out),
    .PE_wrapper290_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper290_U0_fifo_w_out_V_V_din_pass_0_out),
    .fifo_w_PE_11_9_V_V_full_n_pass_0(fifo_w_PE_11_9_V_V_full_n_pass_0_in),
    .PE_wrapper290_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper290_U0_fifo_w_out_V_V_write_pass_0_out),
    .PE_wrapper253_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper253_U0_fifo_cin_out_V_V_din_pass_0_in),
    .fifo_cin_PE_9_7_V_V_full_n_pass_0(fifo_cin_PE_9_7_V_V_full_n_pass_0_out),
    .PE_wrapper253_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper253_U0_fifo_cin_out_V_V_write_pass_0_in),
    .PE_wrapper289_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper289_U0_fifo_cin_out_V_V_din_pass_0_out),
    .fifo_cin_PE_12_7_V_V_full_n_pass_0(fifo_cin_PE_12_7_V_V_full_n_pass_0_in),
    .PE_wrapper289_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper289_U0_fifo_cin_out_V_V_write_pass_0_out),
    .cout_drain_IO_L1_out_wrapper482_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper482_U0_fifo_cout_drain_out_V_V_din_pass_0_in),
    .fifo_cout_drain_cout_drain_IO_L1_out_7_12_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_7_12_V_V_full_n_pass_0_out),
    .cout_drain_IO_L1_out_wrapper482_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper482_U0_fifo_cout_drain_out_V_V_write_pass_0_in),
    .PE_wrapper276_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper276_U0_fifo_w_out_V_V_din_pass_0_in),
    .fifo_w_PE_10_7_V_V_full_n_pass_0(fifo_w_PE_10_7_V_V_full_n_pass_0_out),
    .PE_wrapper276_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper276_U0_fifo_w_out_V_V_write_pass_0_in),
    .PE_wrapper264_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper264_U0_fifo_cout_drain_out_V_din_pass_0_out),
    .fifo_cout_drain_PE_9_6_V_full_n_pass_0(fifo_cout_drain_PE_9_6_V_full_n_pass_0_in),
    .PE_wrapper264_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper264_U0_fifo_cout_drain_out_V_write_pass_0_out),
    .PE_wrapper278_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper278_U0_fifo_w_out_V_V_din_pass_0_out),
    .fifo_w_PE_10_9_V_V_full_n_pass_0(fifo_w_PE_10_9_V_V_full_n_pass_0_in),
    .PE_wrapper278_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper278_U0_fifo_w_out_V_V_write_pass_0_out),
    .PE_wrapper290_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper290_U0_fifo_cin_out_V_V_din_pass_0_out),
    .fifo_cin_PE_12_8_V_V_full_n_pass_0(fifo_cin_PE_12_8_V_V_full_n_pass_0_in),
    .PE_wrapper290_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper290_U0_fifo_cin_out_V_V_write_pass_0_out),
    .cout_drain_IO_L1_out_wrapper497_U0_fifo_cout_drain_out_V_V_din_pass_1(cout_drain_IO_L1_out_wrapper497_U0_fifo_cout_drain_out_V_V_din_pass_1_in),
    .fifo_cout_drain_cout_drain_IO_L1_out_8_13_V_V_full_n_pass_1(fifo_cout_drain_cout_drain_IO_L1_out_8_13_V_V_full_n_pass_1_out),
    .cout_drain_IO_L1_out_wrapper497_U0_fifo_cout_drain_out_V_V_write_pass_1(cout_drain_IO_L1_out_wrapper497_U0_fifo_cout_drain_out_V_V_write_pass_1_in),
    .PE_wrapper264_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper264_U0_fifo_cin_out_V_V_din_pass_0_out),
    .fifo_cin_PE_10_6_V_V_full_n_pass_0(fifo_cin_PE_10_6_V_V_full_n_pass_0_in),
    .PE_wrapper264_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper264_U0_fifo_cin_out_V_V_write_pass_0_out),
    .PE_wrapper252_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper252_U0_fifo_cin_out_V_V_din_pass_0_in),
    .fifo_cin_PE_9_6_V_V_full_n_pass_0(fifo_cin_PE_9_6_V_V_full_n_pass_0_out),
    .PE_wrapper252_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper252_U0_fifo_cin_out_V_V_write_pass_0_in),
    .PE_wrapper302_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper302_U0_fifo_cout_drain_out_V_din_pass_0_in),
    .fifo_cout_drain_PE_12_8_V_full_n_pass_0(fifo_cout_drain_PE_12_8_V_full_n_pass_0_out),
    .PE_wrapper302_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper302_U0_fifo_cout_drain_out_V_write_pass_0_in),
    .PE_wrapper266_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper266_U0_fifo_w_out_V_V_din_pass_0_out),
    .fifo_w_PE_9_9_V_V_full_n_pass_0(fifo_w_PE_9_9_V_V_full_n_pass_0_in),
    .PE_wrapper266_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper266_U0_fifo_w_out_V_V_write_pass_0_out),
    .cout_drain_IO_L1_out_wrapper501_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper501_U0_fifo_cout_drain_out_V_V_din_pass_0_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_8_9_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_8_9_V_V_full_n_pass_0_in),
    .cout_drain_IO_L1_out_wrapper501_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper501_U0_fifo_cout_drain_out_V_V_write_pass_0_out),
    .PE_wrapper263_U0_fifo_w_out_V_V_din_pass_1(PE_wrapper263_U0_fifo_w_out_V_V_din_pass_1_in),
    .fifo_w_PE_9_6_V_V_full_n_pass_1(fifo_w_PE_9_6_V_V_full_n_pass_1_out),
    .PE_wrapper263_U0_fifo_w_out_V_V_write_pass_1(PE_wrapper263_U0_fifo_w_out_V_V_write_pass_1_in),
    .cout_drain_IO_L1_out_wrapper485_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper485_U0_fifo_cout_drain_out_V_V_din_pass_0_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_7_9_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_7_9_V_V_full_n_pass_0_in),
    .cout_drain_IO_L1_out_wrapper485_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper485_U0_fifo_cout_drain_out_V_V_write_pass_0_out),
    .PE_wrapper254_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper254_U0_fifo_cin_out_V_V_din_pass_0_in),
    .fifo_cin_PE_9_8_V_V_full_n_pass_0(fifo_cin_PE_9_8_V_V_full_n_pass_0_out),
    .PE_wrapper254_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper254_U0_fifo_cin_out_V_V_write_pass_0_in),
    .PE_wrapper288_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper288_U0_fifo_w_out_V_V_din_pass_0_in),
    .fifo_w_PE_11_7_V_V_full_n_pass_0(fifo_w_PE_11_7_V_V_full_n_pass_0_out),
    .PE_wrapper288_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper288_U0_fifo_w_out_V_V_write_pass_0_in),
    .ap_clk(ap_clk),
    .ap_start_Boundary_X2Y10_To_X4Y10(ap_start_Boundary_X2Y10_To_X4Y10_in),
    .ap_rst_n_Boundary_X2Y10_To_X4Y10(ap_rst_n_Boundary_X2Y10_To_X4Y10_in),
    .ap_done_Boundary_X2Y10_To_X4Y10(ap_done_Boundary_X2Y10_To_X4Y10_out),
    .ap_start_Boundary_X2Y12_To_X4Y12(ap_start_Boundary_X2Y12_To_X4Y12_out),
    .ap_rst_n_Boundary_X2Y12_To_X4Y12(ap_rst_n_Boundary_X2Y12_To_X4Y12_out),
    .ap_done_Boundary_X2Y12_To_X4Y12(ap_done_Boundary_X2Y12_To_X4Y12_in)
  );


  (* keep_hierarchy = "yes" *) CR_X0Y12_To_CR_X1Y13_ctrl CR_X0Y12_To_CR_X1Y13_ctrl_U0 (
    .PE_wrapper304_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper304_U0_fifo_cin_out_V_V_din_pass_0_in),
    .PE_wrapper304_U0_fifo_cin_out_V_V_din_pass_1(PE_wrapper304_U0_fifo_cin_out_V_V_din_pass_1_out),
    .fifo_cin_PE_13_10_V_V_full_n_pass_0(fifo_cin_PE_13_10_V_V_full_n_pass_0_out),
    .fifo_cin_PE_13_10_V_V_full_n_pass_1(fifo_cin_PE_13_10_V_V_full_n_pass_1_in),
    .PE_wrapper304_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper304_U0_fifo_cin_out_V_V_write_pass_0_in),
    .PE_wrapper304_U0_fifo_cin_out_V_V_write_pass_1(PE_wrapper304_U0_fifo_cin_out_V_V_write_pass_1_out),
    .PE_wrapper305_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper305_U0_fifo_cin_out_V_V_din_pass_0_in),
    .PE_wrapper305_U0_fifo_cin_out_V_V_din_pass_1(PE_wrapper305_U0_fifo_cin_out_V_V_din_pass_1_out),
    .fifo_cin_PE_13_11_V_V_full_n_pass_0(fifo_cin_PE_13_11_V_V_full_n_pass_0_out),
    .fifo_cin_PE_13_11_V_V_full_n_pass_1(fifo_cin_PE_13_11_V_V_full_n_pass_1_in),
    .PE_wrapper305_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper305_U0_fifo_cin_out_V_V_write_pass_0_in),
    .PE_wrapper305_U0_fifo_cin_out_V_V_write_pass_1(PE_wrapper305_U0_fifo_cin_out_V_V_write_pass_1_out),
    .cout_drain_IO_L1_out_wrapper513_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper513_U0_fifo_cout_drain_out_V_V_din_pass_0_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_9_13_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_9_13_V_V_full_n_pass_0_in),
    .cout_drain_IO_L1_out_wrapper513_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper513_U0_fifo_cout_drain_out_V_V_write_pass_0_out),
    .PE_wrapper303_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper303_U0_fifo_cin_out_V_V_din_pass_0_in),
    .fifo_cin_PE_13_9_V_V_full_n_pass_0(fifo_cin_PE_13_9_V_V_full_n_pass_0_out),
    .PE_wrapper303_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper303_U0_fifo_cin_out_V_V_write_pass_0_in),
    .PE_wrapper327_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper327_U0_fifo_w_out_V_V_din_pass_0_out),
    .fifo_w_PE_14_10_V_V_full_n_pass_0(fifo_w_PE_14_10_V_V_full_n_pass_0_in),
    .PE_wrapper327_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper327_U0_fifo_w_out_V_V_write_pass_0_out),
    .cout_drain_IO_L1_out_wrapper497_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper497_U0_fifo_cout_drain_out_V_V_din_pass_0_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_8_13_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_8_13_V_V_full_n_pass_0_in),
    .cout_drain_IO_L1_out_wrapper497_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper497_U0_fifo_cout_drain_out_V_V_write_pass_0_out),
    .PE_wrapper325_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper325_U0_fifo_w_out_V_V_din_pass_0_in),
    .fifo_w_PE_14_8_V_V_full_n_pass_0(fifo_w_PE_14_8_V_V_full_n_pass_0_out),
    .PE_wrapper325_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper325_U0_fifo_w_out_V_V_write_pass_0_in),
    .PE_wrapper315_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper315_U0_fifo_w_out_V_V_din_pass_0_out),
    .fifo_w_PE_13_10_V_V_full_n_pass_0(fifo_w_PE_13_10_V_V_full_n_pass_0_in),
    .PE_wrapper315_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper315_U0_fifo_w_out_V_V_write_pass_0_out),
    .PE_wrapper302_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper302_U0_fifo_cin_out_V_V_din_pass_0_in),
    .fifo_cin_PE_13_8_V_V_full_n_pass_0(fifo_cin_PE_13_8_V_V_full_n_pass_0_out),
    .PE_wrapper302_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper302_U0_fifo_cin_out_V_V_write_pass_0_in),
    .PE_wrapper337_U0_fifo_w_out_V_V_din_pass_1(PE_wrapper337_U0_fifo_w_out_V_V_din_pass_1_in),
    .fifo_w_PE_15_8_V_V_full_n_pass_1(fifo_w_PE_15_8_V_V_full_n_pass_1_out),
    .PE_wrapper337_U0_fifo_w_out_V_V_write_pass_1(PE_wrapper337_U0_fifo_w_out_V_V_write_pass_1_in),
    .PE_wrapper313_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper313_U0_fifo_w_out_V_V_din_pass_0_in),
    .fifo_w_PE_13_8_V_V_full_n_pass_0(fifo_w_PE_13_8_V_V_full_n_pass_0_out),
    .PE_wrapper313_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper313_U0_fifo_w_out_V_V_write_pass_0_in),
    .PE_wrapper339_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper339_U0_fifo_w_out_V_V_din_pass_0_out),
    .fifo_w_PE_15_10_V_V_full_n_pass_0(fifo_w_PE_15_10_V_V_full_n_pass_0_in),
    .PE_wrapper339_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper339_U0_fifo_w_out_V_V_write_pass_0_out),
    .ap_clk(ap_clk),
    .ap_start_Boundary_X0Y12_To_X2Y12(ap_start_Boundary_X0Y12_To_X2Y12_in),
    .ap_rst_n_Boundary_X0Y12_To_X2Y12(ap_rst_n_Boundary_X0Y12_To_X2Y12_in),
    .ap_done_Boundary_X0Y12_To_X2Y12(ap_done_Boundary_X0Y12_To_X2Y12_out),
    .ap_start_Boundary_X0Y14_To_X2Y14(ap_start_Boundary_X0Y14_To_X2Y14_out),
    .ap_rst_n_Boundary_X0Y14_To_X2Y14(ap_rst_n_Boundary_X0Y14_To_X2Y14_out),
    .ap_done_Boundary_X0Y14_To_X2Y14(ap_done_Boundary_X0Y14_To_X2Y14_in)
  );


  (* keep_hierarchy = "yes" *) CR_X0Y14_To_CR_X1Y15_ctrl CR_X0Y14_To_CR_X1Y15_ctrl_U0 (
    .PE_wrapper304_U0_fifo_cin_out_V_V_din_pass_1(PE_wrapper304_U0_fifo_cin_out_V_V_din_pass_1_in),
    .fifo_cin_PE_13_10_V_V_full_n_pass_1(fifo_cin_PE_13_10_V_V_full_n_pass_1_out),
    .PE_wrapper304_U0_fifo_cin_out_V_V_write_pass_1(PE_wrapper304_U0_fifo_cin_out_V_V_write_pass_1_in),
    .PE_wrapper327_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper327_U0_fifo_w_out_V_V_din_pass_0_in),
    .fifo_w_PE_14_10_V_V_full_n_pass_0(fifo_w_PE_14_10_V_V_full_n_pass_0_out),
    .PE_wrapper327_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper327_U0_fifo_w_out_V_V_write_pass_0_in),
    .PE_wrapper315_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper315_U0_fifo_w_out_V_V_din_pass_0_in),
    .fifo_w_PE_13_10_V_V_full_n_pass_0(fifo_w_PE_13_10_V_V_full_n_pass_0_out),
    .PE_wrapper315_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper315_U0_fifo_w_out_V_V_write_pass_0_in),
    .cout_drain_IO_L1_out_wrapper529_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper529_U0_fifo_cout_drain_out_V_V_din_pass_0_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_10_13_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_10_13_V_V_full_n_pass_0_in),
    .cout_drain_IO_L1_out_wrapper529_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper529_U0_fifo_cout_drain_out_V_V_write_pass_0_out),
    .PE_wrapper305_U0_fifo_cin_out_V_V_din_pass_1(PE_wrapper305_U0_fifo_cin_out_V_V_din_pass_1_in),
    .fifo_cin_PE_13_11_V_V_full_n_pass_1(fifo_cin_PE_13_11_V_V_full_n_pass_1_out),
    .PE_wrapper305_U0_fifo_cin_out_V_V_write_pass_1(PE_wrapper305_U0_fifo_cin_out_V_V_write_pass_1_in),
    .PE_wrapper339_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper339_U0_fifo_w_out_V_V_din_pass_0_in),
    .fifo_w_PE_15_10_V_V_full_n_pass_0(fifo_w_PE_15_10_V_V_full_n_pass_0_out),
    .PE_wrapper339_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper339_U0_fifo_w_out_V_V_write_pass_0_in),
    .cout_drain_IO_L1_out_wrapper544_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper544_U0_fifo_cout_drain_out_V_V_din_pass_0_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_11_13_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_11_13_V_V_full_n_pass_0_in),
    .cout_drain_IO_L1_out_wrapper544_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper544_U0_fifo_cout_drain_out_V_V_write_pass_0_out),
    .ap_clk(ap_clk),
    .ap_start_Boundary_X0Y14_To_X2Y14(ap_start_Boundary_X0Y14_To_X2Y14_in),
    .ap_rst_n_Boundary_X0Y14_To_X2Y14(ap_rst_n_Boundary_X0Y14_To_X2Y14_in),
    .ap_done_Boundary_X0Y14_To_X2Y14(ap_done_Boundary_X0Y14_To_X2Y14_out)
  );


  (* keep_hierarchy = "yes" *) CR_X2Y12_To_CR_X3Y13_ctrl CR_X2Y12_To_CR_X3Y13_ctrl_U0 (
    .cout_drain_IO_L1_out_wrapper497_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper497_U0_fifo_cout_drain_out_V_V_din_pass_0_in),
    .cout_drain_IO_L1_out_wrapper497_U0_fifo_cout_drain_out_V_V_din_pass_1(cout_drain_IO_L1_out_wrapper497_U0_fifo_cout_drain_out_V_V_din_pass_1_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_8_13_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_8_13_V_V_full_n_pass_0_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_8_13_V_V_full_n_pass_1(fifo_cout_drain_cout_drain_IO_L1_out_8_13_V_V_full_n_pass_1_in),
    .cout_drain_IO_L1_out_wrapper497_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper497_U0_fifo_cout_drain_out_V_V_write_pass_0_in),
    .cout_drain_IO_L1_out_wrapper497_U0_fifo_cout_drain_out_V_V_write_pass_1(cout_drain_IO_L1_out_wrapper497_U0_fifo_cout_drain_out_V_V_write_pass_1_out),
    .PE_wrapper278_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper278_U0_fifo_w_out_V_V_din_pass_0_in),
    .PE_wrapper278_U0_fifo_w_out_V_V_din_pass_1(PE_wrapper278_U0_fifo_w_out_V_V_din_pass_1_out),
    .fifo_w_PE_10_9_V_V_full_n_pass_0(fifo_w_PE_10_9_V_V_full_n_pass_0_out),
    .fifo_w_PE_10_9_V_V_full_n_pass_1(fifo_w_PE_10_9_V_V_full_n_pass_1_in),
    .PE_wrapper278_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper278_U0_fifo_w_out_V_V_write_pass_0_in),
    .PE_wrapper278_U0_fifo_w_out_V_V_write_pass_1(PE_wrapper278_U0_fifo_w_out_V_V_write_pass_1_out),
    .PE_wrapper290_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper290_U0_fifo_w_out_V_V_din_pass_0_in),
    .fifo_w_PE_11_9_V_V_full_n_pass_0(fifo_w_PE_11_9_V_V_full_n_pass_0_out),
    .PE_wrapper290_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper290_U0_fifo_w_out_V_V_write_pass_0_in),
    .PE_wrapper304_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper304_U0_fifo_cin_out_V_V_din_pass_0_out),
    .fifo_cin_PE_13_10_V_V_full_n_pass_0(fifo_cin_PE_13_10_V_V_full_n_pass_0_in),
    .PE_wrapper304_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper304_U0_fifo_cin_out_V_V_write_pass_0_out),
    .PE_wrapper279_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper279_U0_fifo_cin_out_V_V_din_pass_0_in),
    .fifo_cin_PE_11_9_V_V_full_n_pass_0(fifo_cin_PE_11_9_V_V_full_n_pass_0_out),
    .PE_wrapper279_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper279_U0_fifo_cin_out_V_V_write_pass_0_in),
    .PE_wrapper267_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper267_U0_fifo_cin_out_V_V_din_pass_0_out),
    .fifo_cin_PE_10_9_V_V_full_n_pass_0(fifo_cin_PE_10_9_V_V_full_n_pass_0_in),
    .PE_wrapper267_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper267_U0_fifo_cin_out_V_V_write_pass_0_out),
    .PE_wrapper269_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper269_U0_fifo_cout_drain_out_V_din_pass_0_in),
    .fifo_cout_drain_PE_9_11_V_full_n_pass_0(fifo_cout_drain_PE_9_11_V_full_n_pass_0_out),
    .PE_wrapper269_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper269_U0_fifo_cout_drain_out_V_write_pass_0_in),
    .cout_drain_IO_L1_out_wrapper513_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper513_U0_fifo_cout_drain_out_V_V_din_pass_0_in),
    .fifo_cout_drain_cout_drain_IO_L1_out_9_13_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_9_13_V_V_full_n_pass_0_out),
    .cout_drain_IO_L1_out_wrapper513_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper513_U0_fifo_cout_drain_out_V_V_write_pass_0_in),
    .PE_wrapper292_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper292_U0_fifo_w_out_V_V_din_pass_0_in),
    .fifo_w_PE_11_11_V_V_full_n_pass_0(fifo_w_PE_11_11_V_V_full_n_pass_0_out),
    .PE_wrapper292_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper292_U0_fifo_w_out_V_V_write_pass_0_in),
    .PE_wrapper281_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper281_U0_fifo_cout_drain_out_V_din_pass_0_in),
    .fifo_cout_drain_PE_10_11_V_full_n_pass_0(fifo_cout_drain_PE_10_11_V_full_n_pass_0_out),
    .PE_wrapper281_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper281_U0_fifo_cout_drain_out_V_write_pass_0_in),
    .PE_wrapper280_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper280_U0_fifo_cout_drain_out_V_din_pass_0_in),
    .fifo_cout_drain_PE_10_10_V_full_n_pass_0(fifo_cout_drain_PE_10_10_V_full_n_pass_0_out),
    .PE_wrapper280_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper280_U0_fifo_cout_drain_out_V_write_pass_0_in),
    .PE_wrapper281_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper281_U0_fifo_cin_out_V_V_din_pass_0_in),
    .fifo_cin_PE_11_11_V_V_full_n_pass_0(fifo_cin_PE_11_11_V_V_full_n_pass_0_out),
    .PE_wrapper281_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper281_U0_fifo_cin_out_V_V_write_pass_0_in),
    .PE_wrapper302_U0_fifo_w_out_V_V_din_pass_1(PE_wrapper302_U0_fifo_w_out_V_V_din_pass_1_in),
    .fifo_w_PE_12_9_V_V_full_n_pass_1(fifo_w_PE_12_9_V_V_full_n_pass_1_out),
    .PE_wrapper302_U0_fifo_w_out_V_V_write_pass_1(PE_wrapper302_U0_fifo_w_out_V_V_write_pass_1_in),
    .PE_wrapper291_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper291_U0_fifo_w_out_V_V_din_pass_0_out),
    .fifo_w_PE_11_10_V_V_full_n_pass_0(fifo_w_PE_11_10_V_V_full_n_pass_0_in),
    .PE_wrapper291_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper291_U0_fifo_w_out_V_V_write_pass_0_out),
    .PE_wrapper255_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper255_U0_fifo_cin_out_V_V_din_pass_0_in),
    .fifo_cin_PE_9_9_V_V_full_n_pass_0(fifo_cin_PE_9_9_V_V_full_n_pass_0_out),
    .PE_wrapper255_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper255_U0_fifo_cin_out_V_V_write_pass_0_in),
    .PE_wrapper292_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper292_U0_fifo_cin_out_V_V_din_pass_0_in),
    .fifo_cin_PE_12_10_V_V_full_n_pass_0(fifo_cin_PE_12_10_V_V_full_n_pass_0_out),
    .PE_wrapper292_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper292_U0_fifo_cin_out_V_V_write_pass_0_in),
    .cout_drain_IO_L1_out_wrapper517_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper517_U0_fifo_cout_drain_out_V_V_din_pass_0_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_9_9_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_9_9_V_V_full_n_pass_0_in),
    .cout_drain_IO_L1_out_wrapper517_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper517_U0_fifo_cout_drain_out_V_V_write_pass_0_out),
    .PE_wrapper268_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper268_U0_fifo_cout_drain_out_V_din_pass_0_in),
    .fifo_cout_drain_PE_9_10_V_full_n_pass_0(fifo_cout_drain_PE_9_10_V_full_n_pass_0_out),
    .PE_wrapper268_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper268_U0_fifo_cout_drain_out_V_write_pass_0_in),
    .PE_wrapper266_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper266_U0_fifo_w_out_V_V_din_pass_0_in),
    .fifo_w_PE_9_9_V_V_full_n_pass_0(fifo_w_PE_9_9_V_V_full_n_pass_0_out),
    .PE_wrapper266_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper266_U0_fifo_w_out_V_V_write_pass_0_in),
    .cout_drain_IO_L1_out_wrapper529_U0_fifo_cout_drain_out_V_V_din_pass_1(cout_drain_IO_L1_out_wrapper529_U0_fifo_cout_drain_out_V_V_din_pass_1_in),
    .fifo_cout_drain_cout_drain_IO_L1_out_10_13_V_V_full_n_pass_1(fifo_cout_drain_cout_drain_IO_L1_out_10_13_V_V_full_n_pass_1_out),
    .cout_drain_IO_L1_out_wrapper529_U0_fifo_cout_drain_out_V_V_write_pass_1(cout_drain_IO_L1_out_wrapper529_U0_fifo_cout_drain_out_V_V_write_pass_1_in),
    .cout_drain_IO_L1_out_wrapper533_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper533_U0_fifo_cout_drain_out_V_V_din_pass_0_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_10_9_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_10_9_V_V_full_n_pass_0_in),
    .cout_drain_IO_L1_out_wrapper533_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper533_U0_fifo_cout_drain_out_V_V_write_pass_0_out),
    .PE_wrapper267_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper267_U0_fifo_w_out_V_V_din_pass_0_out),
    .fifo_w_PE_9_10_V_V_full_n_pass_0(fifo_w_PE_9_10_V_V_full_n_pass_0_in),
    .PE_wrapper267_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper267_U0_fifo_w_out_V_V_write_pass_0_out),
    .PE_wrapper305_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper305_U0_fifo_cin_out_V_V_din_pass_0_out),
    .fifo_cin_PE_13_11_V_V_full_n_pass_0(fifo_cin_PE_13_11_V_V_full_n_pass_0_in),
    .PE_wrapper305_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper305_U0_fifo_cin_out_V_V_write_pass_0_out),
    .PE_wrapper292_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper292_U0_fifo_cout_drain_out_V_din_pass_0_in),
    .fifo_cout_drain_PE_11_10_V_full_n_pass_0(fifo_cout_drain_PE_11_10_V_full_n_pass_0_out),
    .PE_wrapper292_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper292_U0_fifo_cout_drain_out_V_write_pass_0_in),
    .cout_drain_IO_L1_out_wrapper548_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper548_U0_fifo_cout_drain_out_V_V_din_pass_0_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_11_9_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_11_9_V_V_full_n_pass_0_in),
    .cout_drain_IO_L1_out_wrapper548_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper548_U0_fifo_cout_drain_out_V_V_write_pass_0_out),
    .PE_wrapper279_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper279_U0_fifo_cout_drain_out_V_din_pass_0_in),
    .fifo_cout_drain_PE_10_9_V_full_n_pass_0(fifo_cout_drain_PE_10_9_V_full_n_pass_0_out),
    .PE_wrapper279_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper279_U0_fifo_cout_drain_out_V_write_pass_0_in),
    .PE_wrapper303_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper303_U0_fifo_cin_out_V_V_din_pass_0_out),
    .fifo_cin_PE_13_9_V_V_full_n_pass_0(fifo_cin_PE_13_9_V_V_full_n_pass_0_in),
    .PE_wrapper303_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper303_U0_fifo_cin_out_V_V_write_pass_0_out),
    .cout_drain_IO_L1_out_wrapper544_U0_fifo_cout_drain_out_V_V_din_pass_1(cout_drain_IO_L1_out_wrapper544_U0_fifo_cout_drain_out_V_V_din_pass_1_in),
    .fifo_cout_drain_cout_drain_IO_L1_out_11_13_V_V_full_n_pass_1(fifo_cout_drain_cout_drain_IO_L1_out_11_13_V_V_full_n_pass_1_out),
    .cout_drain_IO_L1_out_wrapper544_U0_fifo_cout_drain_out_V_V_write_pass_1(cout_drain_IO_L1_out_wrapper544_U0_fifo_cout_drain_out_V_V_write_pass_1_in),
    .ap_clk(ap_clk),
    .ap_start_Boundary_X2Y12_To_X4Y12(ap_start_Boundary_X2Y12_To_X4Y12_in),
    .ap_rst_n_Boundary_X2Y12_To_X4Y12(ap_rst_n_Boundary_X2Y12_To_X4Y12_in),
    .ap_done_Boundary_X2Y12_To_X4Y12(ap_done_Boundary_X2Y12_To_X4Y12_out),
    .ap_start_Boundary_X2Y14_To_X4Y14(ap_start_Boundary_X2Y14_To_X4Y14_out),
    .ap_rst_n_Boundary_X2Y14_To_X4Y14(ap_rst_n_Boundary_X2Y14_To_X4Y14_out),
    .ap_done_Boundary_X2Y14_To_X4Y14(ap_done_Boundary_X2Y14_To_X4Y14_in)
  );


  (* keep_hierarchy = "yes" *) CR_X2Y14_To_CR_X3Y15_ctrl CR_X2Y14_To_CR_X3Y15_ctrl_U0 (
    .cout_drain_IO_L1_out_wrapper529_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper529_U0_fifo_cout_drain_out_V_V_din_pass_0_in),
    .cout_drain_IO_L1_out_wrapper529_U0_fifo_cout_drain_out_V_V_din_pass_1(cout_drain_IO_L1_out_wrapper529_U0_fifo_cout_drain_out_V_V_din_pass_1_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_10_13_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_10_13_V_V_full_n_pass_0_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_10_13_V_V_full_n_pass_1(fifo_cout_drain_cout_drain_IO_L1_out_10_13_V_V_full_n_pass_1_in),
    .cout_drain_IO_L1_out_wrapper529_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper529_U0_fifo_cout_drain_out_V_V_write_pass_0_in),
    .cout_drain_IO_L1_out_wrapper529_U0_fifo_cout_drain_out_V_V_write_pass_1(cout_drain_IO_L1_out_wrapper529_U0_fifo_cout_drain_out_V_V_write_pass_1_out),
    .cout_drain_IO_L1_out_wrapper544_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper544_U0_fifo_cout_drain_out_V_V_din_pass_0_in),
    .cout_drain_IO_L1_out_wrapper544_U0_fifo_cout_drain_out_V_V_din_pass_1(cout_drain_IO_L1_out_wrapper544_U0_fifo_cout_drain_out_V_V_din_pass_1_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_11_13_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_11_13_V_V_full_n_pass_0_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_11_13_V_V_full_n_pass_1(fifo_cout_drain_cout_drain_IO_L1_out_11_13_V_V_full_n_pass_1_in),
    .cout_drain_IO_L1_out_wrapper544_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper544_U0_fifo_cout_drain_out_V_V_write_pass_0_in),
    .cout_drain_IO_L1_out_wrapper544_U0_fifo_cout_drain_out_V_V_write_pass_1(cout_drain_IO_L1_out_wrapper544_U0_fifo_cout_drain_out_V_V_write_pass_1_out),
    .PE_wrapper279_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper279_U0_fifo_cin_out_V_V_din_pass_0_out),
    .fifo_cin_PE_11_9_V_V_full_n_pass_0(fifo_cin_PE_11_9_V_V_full_n_pass_0_in),
    .PE_wrapper279_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper279_U0_fifo_cin_out_V_V_write_pass_0_out),
    .PE_wrapper269_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper269_U0_fifo_cout_drain_out_V_din_pass_0_out),
    .fifo_cout_drain_PE_9_11_V_full_n_pass_0(fifo_cout_drain_PE_9_11_V_full_n_pass_0_in),
    .PE_wrapper269_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper269_U0_fifo_cout_drain_out_V_write_pass_0_out),
    .PE_wrapper267_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper267_U0_fifo_cin_out_V_V_din_pass_0_in),
    .fifo_cin_PE_10_9_V_V_full_n_pass_0(fifo_cin_PE_10_9_V_V_full_n_pass_0_out),
    .PE_wrapper267_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper267_U0_fifo_cin_out_V_V_write_pass_0_in),
    .PE_wrapper292_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper292_U0_fifo_w_out_V_V_din_pass_0_out),
    .fifo_w_PE_11_11_V_V_full_n_pass_0(fifo_w_PE_11_11_V_V_full_n_pass_0_in),
    .PE_wrapper292_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper292_U0_fifo_w_out_V_V_write_pass_0_out),
    .PE_wrapper281_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper281_U0_fifo_cout_drain_out_V_din_pass_0_out),
    .fifo_cout_drain_PE_10_11_V_full_n_pass_0(fifo_cout_drain_PE_10_11_V_full_n_pass_0_in),
    .PE_wrapper281_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper281_U0_fifo_cout_drain_out_V_write_pass_0_out),
    .PE_wrapper280_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper280_U0_fifo_cout_drain_out_V_din_pass_0_out),
    .fifo_cout_drain_PE_10_10_V_full_n_pass_0(fifo_cout_drain_PE_10_10_V_full_n_pass_0_in),
    .PE_wrapper280_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper280_U0_fifo_cout_drain_out_V_write_pass_0_out),
    .PE_wrapper278_U0_fifo_w_out_V_V_din_pass_1(PE_wrapper278_U0_fifo_w_out_V_V_din_pass_1_in),
    .fifo_w_PE_10_9_V_V_full_n_pass_1(fifo_w_PE_10_9_V_V_full_n_pass_1_out),
    .PE_wrapper278_U0_fifo_w_out_V_V_write_pass_1(PE_wrapper278_U0_fifo_w_out_V_V_write_pass_1_in),
    .PE_wrapper281_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper281_U0_fifo_cin_out_V_V_din_pass_0_out),
    .fifo_cin_PE_11_11_V_V_full_n_pass_0(fifo_cin_PE_11_11_V_V_full_n_pass_0_in),
    .PE_wrapper281_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper281_U0_fifo_cin_out_V_V_write_pass_0_out),
    .PE_wrapper256_U0_fifo_cin_out_V_V_din_pass_1(PE_wrapper256_U0_fifo_cin_out_V_V_din_pass_1_in),
    .fifo_cin_PE_9_10_V_V_full_n_pass_1(fifo_cin_PE_9_10_V_V_full_n_pass_1_out),
    .PE_wrapper256_U0_fifo_cin_out_V_V_write_pass_1(PE_wrapper256_U0_fifo_cin_out_V_V_write_pass_1_in),
    .PE_wrapper291_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper291_U0_fifo_w_out_V_V_din_pass_0_in),
    .fifo_w_PE_11_10_V_V_full_n_pass_0(fifo_w_PE_11_10_V_V_full_n_pass_0_out),
    .PE_wrapper291_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper291_U0_fifo_w_out_V_V_write_pass_0_in),
    .PE_wrapper292_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper292_U0_fifo_cin_out_V_V_din_pass_0_out),
    .fifo_cin_PE_12_10_V_V_full_n_pass_0(fifo_cin_PE_12_10_V_V_full_n_pass_0_in),
    .PE_wrapper292_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper292_U0_fifo_cin_out_V_V_write_pass_0_out),
    .PE_wrapper268_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper268_U0_fifo_cout_drain_out_V_din_pass_0_out),
    .fifo_cout_drain_PE_9_10_V_full_n_pass_0(fifo_cout_drain_PE_9_10_V_full_n_pass_0_in),
    .PE_wrapper268_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper268_U0_fifo_cout_drain_out_V_write_pass_0_out),
    .PE_wrapper257_U0_fifo_cin_out_V_V_din_pass_1(PE_wrapper257_U0_fifo_cin_out_V_V_din_pass_1_in),
    .fifo_cin_PE_9_11_V_V_full_n_pass_1(fifo_cin_PE_9_11_V_V_full_n_pass_1_out),
    .PE_wrapper257_U0_fifo_cin_out_V_V_write_pass_1(PE_wrapper257_U0_fifo_cin_out_V_V_write_pass_1_in),
    .PE_wrapper267_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper267_U0_fifo_w_out_V_V_din_pass_0_in),
    .fifo_w_PE_9_10_V_V_full_n_pass_0(fifo_w_PE_9_10_V_V_full_n_pass_0_out),
    .PE_wrapper267_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper267_U0_fifo_w_out_V_V_write_pass_0_in),
    .PE_wrapper292_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper292_U0_fifo_cout_drain_out_V_din_pass_0_out),
    .fifo_cout_drain_PE_11_10_V_full_n_pass_0(fifo_cout_drain_PE_11_10_V_full_n_pass_0_in),
    .PE_wrapper292_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper292_U0_fifo_cout_drain_out_V_write_pass_0_out),
    .PE_wrapper279_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper279_U0_fifo_cout_drain_out_V_din_pass_0_out),
    .fifo_cout_drain_PE_10_9_V_full_n_pass_0(fifo_cout_drain_PE_10_9_V_full_n_pass_0_in),
    .PE_wrapper279_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper279_U0_fifo_cout_drain_out_V_write_pass_0_out),
    .ap_clk(ap_clk),
    .ap_start_Boundary_X2Y14_To_X4Y14(ap_start_Boundary_X2Y14_To_X4Y14_in),
    .ap_rst_n_Boundary_X2Y14_To_X4Y14(ap_rst_n_Boundary_X2Y14_To_X4Y14_in),
    .ap_done_Boundary_X2Y14_To_X4Y14(ap_done_Boundary_X2Y14_To_X4Y14_out)
  );


  (* keep_hierarchy = "yes" *) CR_X4Y2_To_CR_X5Y3_ctrl CR_X4Y2_To_CR_X5Y3_ctrl_U0 (
    .w_IO_L2_in140_U0_fifo_w_out_V_V_din_pass_0(w_IO_L2_in140_U0_fifo_w_out_V_V_din_pass_0_in),
    .w_IO_L2_in140_U0_fifo_w_out_V_V_din_pass_1(w_IO_L2_in140_U0_fifo_w_out_V_V_din_pass_1_out),
    .fifo_w_w_IO_L2_in_6_V_V_full_n_pass_0(fifo_w_w_IO_L2_in_6_V_V_full_n_pass_0_out),
    .fifo_w_w_IO_L2_in_6_V_V_full_n_pass_1(fifo_w_w_IO_L2_in_6_V_V_full_n_pass_1_in),
    .w_IO_L2_in140_U0_fifo_w_out_V_V_write_pass_0(w_IO_L2_in140_U0_fifo_w_out_V_V_write_pass_0_in),
    .w_IO_L2_in140_U0_fifo_w_out_V_V_write_pass_1(w_IO_L2_in140_U0_fifo_w_out_V_V_write_pass_1_out),
    .PE_wrapper210_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper210_U0_fifo_cin_out_V_V_din_pass_0_in),
    .PE_wrapper210_U0_fifo_cin_out_V_V_din_pass_1(PE_wrapper210_U0_fifo_cin_out_V_V_din_pass_1_out),
    .fifo_cin_PE_6_0_V_V_full_n_pass_0(fifo_cin_PE_6_0_V_V_full_n_pass_0_out),
    .fifo_cin_PE_6_0_V_V_full_n_pass_1(fifo_cin_PE_6_0_V_V_full_n_pass_1_in),
    .PE_wrapper210_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper210_U0_fifo_cin_out_V_V_write_pass_0_in),
    .PE_wrapper210_U0_fifo_cin_out_V_V_write_pass_1(PE_wrapper210_U0_fifo_cin_out_V_V_write_pass_1_out),
    .w_IO_L2_in138_U0_fifo_w_local_out_V_V_din_pass_0(w_IO_L2_in138_U0_fifo_w_local_out_V_V_din_pass_0_in),
    .w_IO_L2_in138_U0_fifo_w_local_out_V_V_din_pass_1(w_IO_L2_in138_U0_fifo_w_local_out_V_V_din_pass_1_out),
    .fifo_w_PE_3_0_V_V_full_n_pass_0(fifo_w_PE_3_0_V_V_full_n_pass_0_out),
    .fifo_w_PE_3_0_V_V_full_n_pass_1(fifo_w_PE_3_0_V_V_full_n_pass_1_in),
    .w_IO_L2_in138_U0_fifo_w_local_out_V_V_write_pass_0(w_IO_L2_in138_U0_fifo_w_local_out_V_V_write_pass_0_in),
    .w_IO_L2_in138_U0_fifo_w_local_out_V_V_write_pass_1(w_IO_L2_in138_U0_fifo_w_local_out_V_V_write_pass_1_out),
    .cout_drain_IO_L1_out_wrapper378_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper378_U0_fifo_cout_drain_out_V_V_din_pass_0_in),
    .cout_drain_IO_L1_out_wrapper378_U0_fifo_cout_drain_out_V_V_din_pass_1(cout_drain_IO_L1_out_wrapper378_U0_fifo_cout_drain_out_V_V_din_pass_1_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_0_4_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_0_4_V_V_full_n_pass_0_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_0_4_V_V_full_n_pass_1(fifo_cout_drain_cout_drain_IO_L1_out_0_4_V_V_full_n_pass_1_in),
    .cout_drain_IO_L1_out_wrapper378_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper378_U0_fifo_cout_drain_out_V_V_write_pass_0_in),
    .cout_drain_IO_L1_out_wrapper378_U0_fifo_cout_drain_out_V_V_write_pass_1(cout_drain_IO_L1_out_wrapper378_U0_fifo_cout_drain_out_V_V_write_pass_1_out),
    .PE_wrapper201_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper201_U0_fifo_w_out_V_V_din_pass_0_in),
    .PE_wrapper201_U0_fifo_w_out_V_V_din_pass_1(PE_wrapper201_U0_fifo_w_out_V_V_din_pass_1_out),
    .fifo_w_PE_4_4_V_V_full_n_pass_0(fifo_w_PE_4_4_V_V_full_n_pass_0_out),
    .fifo_w_PE_4_4_V_V_full_n_pass_1(fifo_w_PE_4_4_V_V_full_n_pass_1_in),
    .PE_wrapper201_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper201_U0_fifo_w_out_V_V_write_pass_0_in),
    .PE_wrapper201_U0_fifo_w_out_V_V_write_pass_1(PE_wrapper201_U0_fifo_w_out_V_V_write_pass_1_out),
    .PE_wrapper213_U0_fifo_w_out_V_V_din_pass_1(PE_wrapper213_U0_fifo_w_out_V_V_din_pass_1_in),
    .PE_wrapper213_U0_fifo_w_out_V_V_din_pass_2(PE_wrapper213_U0_fifo_w_out_V_V_din_pass_2_out),
    .fifo_w_PE_5_4_V_V_full_n_pass_1(fifo_w_PE_5_4_V_V_full_n_pass_1_out),
    .fifo_w_PE_5_4_V_V_full_n_pass_2(fifo_w_PE_5_4_V_V_full_n_pass_2_in),
    .PE_wrapper213_U0_fifo_w_out_V_V_write_pass_1(PE_wrapper213_U0_fifo_w_out_V_V_write_pass_1_in),
    .PE_wrapper213_U0_fifo_w_out_V_V_write_pass_2(PE_wrapper213_U0_fifo_w_out_V_V_write_pass_2_out),
    .kernel0_entry12_U0_w_V_out_din_pass_0(kernel0_entry12_U0_w_V_out_din_pass_0_in),
    .kernel0_entry12_U0_w_V_out_din_pass_1(kernel0_entry12_U0_w_V_out_din_pass_1_out),
    .w_V_c_full_n_pass_0(w_V_c_full_n_pass_0_out),
    .w_V_c_full_n_pass_1(w_V_c_full_n_pass_1_in),
    .kernel0_entry12_U0_w_V_out_write_pass_0(kernel0_entry12_U0_w_V_out_write_pass_0_in),
    .kernel0_entry12_U0_w_V_out_write_pass_1(kernel0_entry12_U0_w_V_out_write_pass_1_out),
    .kernel0_entry12_U0_cout_V_out_din_pass_0(kernel0_entry12_U0_cout_V_out_din_pass_0_in),
    .kernel0_entry12_U0_cout_V_out_din_pass_1(kernel0_entry12_U0_cout_V_out_din_pass_1_out),
    .cout_V_c_full_n_pass_0(cout_V_c_full_n_pass_0_out),
    .cout_V_c_full_n_pass_1(cout_V_c_full_n_pass_1_in),
    .kernel0_entry12_U0_cout_V_out_write_pass_0(kernel0_entry12_U0_cout_V_out_write_pass_0_in),
    .kernel0_entry12_U0_cout_V_out_write_pass_1(kernel0_entry12_U0_cout_V_out_write_pass_1_out),
    .PE_wrapper165_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper165_U0_fifo_w_out_V_V_din_pass_0_out),
    .fifo_w_PE_1_4_V_V_full_n_pass_0(fifo_w_PE_1_4_V_V_full_n_pass_0_in),
    .PE_wrapper165_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper165_U0_fifo_w_out_V_V_write_pass_0_out),
    .cin_IO_L2_in127_U0_fifo_cin_out_V_V_din_pass_0(cin_IO_L2_in127_U0_fifo_cin_out_V_V_din_pass_0_out),
    .fifo_cin_cin_IO_L2_in_4_V_V_full_n_pass_0(fifo_cin_cin_IO_L2_in_4_V_V_full_n_pass_0_in),
    .cin_IO_L2_in127_U0_fifo_cin_out_V_V_write_pass_0(cin_IO_L2_in127_U0_fifo_cin_out_V_V_write_pass_0_out),
    .PE_wrapper163_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper163_U0_fifo_w_out_V_V_din_pass_0_in),
    .fifo_w_PE_1_2_V_V_full_n_pass_0(fifo_w_PE_1_2_V_V_full_n_pass_0_out),
    .PE_wrapper163_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper163_U0_fifo_w_out_V_V_write_pass_0_in),
    .PE_wrapper188_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper188_U0_fifo_w_out_V_V_din_pass_0_in),
    .fifo_w_PE_3_3_V_V_full_n_pass_0(fifo_w_PE_3_3_V_V_full_n_pass_0_out),
    .PE_wrapper188_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper188_U0_fifo_w_out_V_V_write_pass_0_in),
    .w_IO_L2_in136_U0_fifo_w_out_V_V_din_pass_0(w_IO_L2_in136_U0_fifo_w_out_V_V_din_pass_0_out),
    .fifo_w_w_IO_L2_in_2_V_V_full_n_pass_0(fifo_w_w_IO_L2_in_2_V_V_full_n_pass_0_in),
    .w_IO_L2_in136_U0_fifo_w_out_V_V_write_pass_0(w_IO_L2_in136_U0_fifo_w_out_V_V_write_pass_0_out),
    .PE_wrapper153_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper153_U0_fifo_w_out_V_V_din_pass_0_out),
    .fifo_w_PE_0_4_V_V_full_n_pass_0(fifo_w_PE_0_4_V_V_full_n_pass_0_in),
    .PE_wrapper153_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper153_U0_fifo_w_out_V_V_write_pass_0_out),
    .PE_wrapper177_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper177_U0_fifo_w_out_V_V_din_pass_0_out),
    .fifo_w_PE_2_4_V_V_full_n_pass_0(fifo_w_PE_2_4_V_V_full_n_pass_0_in),
    .PE_wrapper177_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper177_U0_fifo_w_out_V_V_write_pass_0_out),
    .PE_wrapper151_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper151_U0_fifo_w_out_V_V_din_pass_0_in),
    .fifo_w_PE_0_2_V_V_full_n_pass_0(fifo_w_PE_0_2_V_V_full_n_pass_0_out),
    .PE_wrapper151_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper151_U0_fifo_w_out_V_V_write_pass_0_in),
    .PE_wrapper165_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper165_U0_fifo_cout_drain_out_V_din_pass_0_out),
    .fifo_cout_drain_PE_1_3_V_full_n_pass_0(fifo_cout_drain_PE_1_3_V_full_n_pass_0_in),
    .PE_wrapper165_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper165_U0_fifo_cout_drain_out_V_write_pass_0_out),
    .PE_wrapper150_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper150_U0_fifo_cin_out_V_V_din_pass_0_in),
    .fifo_cin_PE_1_0_V_V_full_n_pass_0(fifo_cin_PE_1_0_V_V_full_n_pass_0_out),
    .PE_wrapper150_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper150_U0_fifo_cin_out_V_V_write_pass_0_in),
    .PE_wrapper153_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper153_U0_fifo_cout_drain_out_V_din_pass_0_out),
    .fifo_cout_drain_PE_0_3_V_full_n_pass_0(fifo_cout_drain_PE_0_3_V_full_n_pass_0_in),
    .PE_wrapper153_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper153_U0_fifo_cout_drain_out_V_write_pass_0_out),
    .PE_wrapper177_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper177_U0_fifo_cout_drain_out_V_din_pass_0_out),
    .fifo_cout_drain_PE_2_3_V_full_n_pass_0(fifo_cout_drain_PE_2_3_V_full_n_pass_0_in),
    .PE_wrapper177_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper177_U0_fifo_cout_drain_out_V_write_pass_0_out),
    .PE_wrapper164_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper164_U0_fifo_cout_drain_out_V_din_pass_0_out),
    .fifo_cout_drain_PE_1_2_V_full_n_pass_0(fifo_cout_drain_PE_1_2_V_full_n_pass_0_in),
    .PE_wrapper164_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper164_U0_fifo_cout_drain_out_V_write_pass_0_out),
    .PE_wrapper189_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper189_U0_fifo_cout_drain_out_V_din_pass_0_out),
    .fifo_cout_drain_PE_3_3_V_full_n_pass_0(fifo_cout_drain_PE_3_3_V_full_n_pass_0_in),
    .PE_wrapper189_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper189_U0_fifo_cout_drain_out_V_write_pass_0_out),
    .PE_wrapper162_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper162_U0_fifo_cin_out_V_V_din_pass_0_out),
    .fifo_cin_PE_2_0_V_V_full_n_pass_0(fifo_cin_PE_2_0_V_V_full_n_pass_0_in),
    .PE_wrapper162_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper162_U0_fifo_cin_out_V_V_write_pass_0_out),
    .w_IO_L3_in_serialize_U0_fifo_w_local_out_V_V_din_pass_0(w_IO_L3_in_serialize_U0_fifo_w_local_out_V_V_din_pass_0_in),
    .fifo_w_w_IO_L3_in_serialize_V_V_full_n_pass_0(fifo_w_w_IO_L3_in_serialize_V_V_full_n_pass_0_out),
    .w_IO_L3_in_serialize_U0_fifo_w_local_out_V_V_write_pass_0(w_IO_L3_in_serialize_U0_fifo_w_local_out_V_V_write_pass_0_in),
    .cin_IO_L2_in125_U0_fifo_cin_out_V_V_din_pass_1(cin_IO_L2_in125_U0_fifo_cin_out_V_V_din_pass_1_in),
    .fifo_cin_cin_IO_L2_in_2_V_V_full_n_pass_1(fifo_cin_cin_IO_L2_in_2_V_V_full_n_pass_1_out),
    .cin_IO_L2_in125_U0_fifo_cin_out_V_V_write_pass_1(cin_IO_L2_in125_U0_fifo_cin_out_V_V_write_pass_1_in),
    .PE_wrapper152_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper152_U0_fifo_cout_drain_out_V_din_pass_0_out),
    .fifo_cout_drain_PE_0_2_V_full_n_pass_0(fifo_cout_drain_PE_0_2_V_full_n_pass_0_in),
    .PE_wrapper152_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper152_U0_fifo_cout_drain_out_V_write_pass_0_out),
    .PE_wrapper189_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper189_U0_fifo_w_out_V_V_din_pass_0_out),
    .fifo_w_PE_3_4_V_V_full_n_pass_0(fifo_w_PE_3_4_V_V_full_n_pass_0_in),
    .PE_wrapper189_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper189_U0_fifo_w_out_V_V_write_pass_0_out),
    .PE_wrapper175_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper175_U0_fifo_w_out_V_V_din_pass_0_in),
    .fifo_w_PE_2_2_V_V_full_n_pass_0(fifo_w_PE_2_2_V_V_full_n_pass_0_out),
    .PE_wrapper175_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper175_U0_fifo_w_out_V_V_write_pass_0_in),
    .PE_wrapper162_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper162_U0_fifo_w_out_V_V_din_pass_0_out),
    .fifo_w_PE_1_1_V_V_full_n_pass_0(fifo_w_PE_1_1_V_V_full_n_pass_0_in),
    .PE_wrapper162_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper162_U0_fifo_w_out_V_V_write_pass_0_out),
    .PE_wrapper189_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper189_U0_fifo_cin_out_V_V_din_pass_0_out),
    .fifo_cin_PE_4_3_V_V_full_n_pass_0(fifo_cin_PE_4_3_V_V_full_n_pass_0_in),
    .PE_wrapper189_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper189_U0_fifo_cin_out_V_V_write_pass_0_out),
    .PE_wrapper176_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper176_U0_fifo_cout_drain_out_V_din_pass_0_out),
    .fifo_cout_drain_PE_2_2_V_full_n_pass_0(fifo_cout_drain_PE_2_2_V_full_n_pass_0_in),
    .PE_wrapper176_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper176_U0_fifo_cout_drain_out_V_write_pass_0_out),
    .PE_wrapper176_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper176_U0_fifo_cin_out_V_V_din_pass_0_out),
    .fifo_cin_PE_3_2_V_V_full_n_pass_0(fifo_cin_PE_3_2_V_V_full_n_pass_0_in),
    .PE_wrapper176_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper176_U0_fifo_cin_out_V_V_write_pass_0_out),
    .PE_wrapper162_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper162_U0_fifo_cout_drain_out_V_din_pass_0_out),
    .fifo_cout_drain_PE_1_0_V_full_n_pass_0(fifo_cout_drain_PE_1_0_V_full_n_pass_0_in),
    .PE_wrapper162_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper162_U0_fifo_cout_drain_out_V_write_pass_0_out),
    .w_IO_L2_in135_U0_fifo_w_local_out_V_V_din_pass_0(w_IO_L2_in135_U0_fifo_w_local_out_V_V_din_pass_0_out),
    .fifo_w_PE_0_0_V_V_full_n_pass_0(fifo_w_PE_0_0_V_V_full_n_pass_0_in),
    .w_IO_L2_in135_U0_fifo_w_local_out_V_V_write_pass_0(w_IO_L2_in135_U0_fifo_w_local_out_V_V_write_pass_0_out),
    .ap_clk(ap_clk),
    .ap_start_Boundary_X4Y2_To_X6Y2(ap_start_Boundary_X4Y2_To_X6Y2_in),
    .ap_rst_n_Boundary_X4Y2_To_X6Y2(ap_rst_n_Boundary_X4Y2_To_X6Y2_in),
    .ap_done_Boundary_X4Y2_To_X6Y2(ap_done_Boundary_X4Y2_To_X6Y2_out),
    .ap_start_Boundary_X4Y4_To_X6Y4(ap_start_Boundary_X4Y4_To_X6Y4_out),
    .ap_rst_n_Boundary_X4Y4_To_X6Y4(ap_rst_n_Boundary_X4Y4_To_X6Y4_out),
    .ap_done_Boundary_X4Y4_To_X6Y4(ap_done_Boundary_X4Y4_To_X6Y4_in)
  );


  (* keep_hierarchy = "yes" *) CR_X6Y0_To_CR_X7Y1_ctrl CR_X6Y0_To_CR_X7Y1_ctrl_U0 (
    .PE_wrapper187_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper187_U0_fifo_w_out_V_V_din_pass_0_in),
    .PE_wrapper187_U0_fifo_w_out_V_V_din_pass_1(PE_wrapper187_U0_fifo_w_out_V_V_din_pass_1_out),
    .fifo_w_PE_3_2_V_V_full_n_pass_0(fifo_w_PE_3_2_V_V_full_n_pass_0_out),
    .fifo_w_PE_3_2_V_V_full_n_pass_1(fifo_w_PE_3_2_V_V_full_n_pass_1_in),
    .PE_wrapper187_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper187_U0_fifo_w_out_V_V_write_pass_0_in),
    .PE_wrapper187_U0_fifo_w_out_V_V_write_pass_1(PE_wrapper187_U0_fifo_w_out_V_V_write_pass_1_out),
    .PE_wrapper163_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper163_U0_fifo_cout_drain_out_V_din_pass_0_in),
    .PE_wrapper163_U0_fifo_cout_drain_out_V_din_pass_1(PE_wrapper163_U0_fifo_cout_drain_out_V_din_pass_1_out),
    .fifo_cout_drain_PE_1_1_V_full_n_pass_0(fifo_cout_drain_PE_1_1_V_full_n_pass_0_out),
    .fifo_cout_drain_PE_1_1_V_full_n_pass_1(fifo_cout_drain_PE_1_1_V_full_n_pass_1_in),
    .PE_wrapper163_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper163_U0_fifo_cout_drain_out_V_write_pass_0_in),
    .PE_wrapper163_U0_fifo_cout_drain_out_V_write_pass_1(PE_wrapper163_U0_fifo_cout_drain_out_V_write_pass_1_out),
    .PE_wrapper175_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper175_U0_fifo_cout_drain_out_V_din_pass_0_in),
    .PE_wrapper175_U0_fifo_cout_drain_out_V_din_pass_1(PE_wrapper175_U0_fifo_cout_drain_out_V_din_pass_1_out),
    .fifo_cout_drain_PE_2_1_V_full_n_pass_0(fifo_cout_drain_PE_2_1_V_full_n_pass_0_out),
    .fifo_cout_drain_PE_2_1_V_full_n_pass_1(fifo_cout_drain_PE_2_1_V_full_n_pass_1_in),
    .PE_wrapper175_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper175_U0_fifo_cout_drain_out_V_write_pass_0_in),
    .PE_wrapper175_U0_fifo_cout_drain_out_V_write_pass_1(PE_wrapper175_U0_fifo_cout_drain_out_V_write_pass_1_out),
    .PE_wrapper187_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper187_U0_fifo_cin_out_V_V_din_pass_0_in),
    .PE_wrapper187_U0_fifo_cin_out_V_V_din_pass_1(PE_wrapper187_U0_fifo_cin_out_V_V_din_pass_1_out),
    .fifo_cin_PE_4_1_V_V_full_n_pass_0(fifo_cin_PE_4_1_V_V_full_n_pass_0_out),
    .fifo_cin_PE_4_1_V_V_full_n_pass_1(fifo_cin_PE_4_1_V_V_full_n_pass_1_in),
    .PE_wrapper187_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper187_U0_fifo_cin_out_V_V_write_pass_0_in),
    .PE_wrapper187_U0_fifo_cin_out_V_V_write_pass_1(PE_wrapper187_U0_fifo_cin_out_V_V_write_pass_1_out),
    .PE_wrapper186_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper186_U0_fifo_cin_out_V_V_din_pass_0_in),
    .PE_wrapper186_U0_fifo_cin_out_V_V_din_pass_1(PE_wrapper186_U0_fifo_cin_out_V_V_din_pass_1_out),
    .fifo_cin_PE_4_0_V_V_full_n_pass_0(fifo_cin_PE_4_0_V_V_full_n_pass_0_out),
    .fifo_cin_PE_4_0_V_V_full_n_pass_1(fifo_cin_PE_4_0_V_V_full_n_pass_1_in),
    .PE_wrapper186_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper186_U0_fifo_cin_out_V_V_write_pass_0_in),
    .PE_wrapper186_U0_fifo_cin_out_V_V_write_pass_1(PE_wrapper186_U0_fifo_cin_out_V_V_write_pass_1_out),
    .PE_wrapper187_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper187_U0_fifo_cout_drain_out_V_din_pass_0_in),
    .PE_wrapper187_U0_fifo_cout_drain_out_V_din_pass_1(PE_wrapper187_U0_fifo_cout_drain_out_V_din_pass_1_out),
    .fifo_cout_drain_PE_3_1_V_full_n_pass_0(fifo_cout_drain_PE_3_1_V_full_n_pass_0_out),
    .fifo_cout_drain_PE_3_1_V_full_n_pass_1(fifo_cout_drain_PE_3_1_V_full_n_pass_1_in),
    .PE_wrapper187_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper187_U0_fifo_cout_drain_out_V_write_pass_0_in),
    .PE_wrapper187_U0_fifo_cout_drain_out_V_write_pass_1(PE_wrapper187_U0_fifo_cout_drain_out_V_write_pass_1_out),
    .w_IO_L2_in137_U0_fifo_w_out_V_V_din_pass_0(w_IO_L2_in137_U0_fifo_w_out_V_V_din_pass_0_in),
    .w_IO_L2_in137_U0_fifo_w_out_V_V_din_pass_1(w_IO_L2_in137_U0_fifo_w_out_V_V_din_pass_1_out),
    .fifo_w_w_IO_L2_in_3_V_V_full_n_pass_0(fifo_w_w_IO_L2_in_3_V_V_full_n_pass_0_out),
    .fifo_w_w_IO_L2_in_3_V_V_full_n_pass_1(fifo_w_w_IO_L2_in_3_V_V_full_n_pass_1_in),
    .w_IO_L2_in137_U0_fifo_w_out_V_V_write_pass_0(w_IO_L2_in137_U0_fifo_w_out_V_V_write_pass_0_in),
    .w_IO_L2_in137_U0_fifo_w_out_V_V_write_pass_1(w_IO_L2_in137_U0_fifo_w_out_V_V_write_pass_1_out),
    .cout_drain_IO_L1_out_wrapper376_U0_fifo_cout_drain_out_V_V_din_pass_1(cout_drain_IO_L1_out_wrapper376_U0_fifo_cout_drain_out_V_V_din_pass_1_in),
    .cout_drain_IO_L1_out_wrapper376_U0_fifo_cout_drain_out_V_V_din_pass_2(cout_drain_IO_L1_out_wrapper376_U0_fifo_cout_drain_out_V_V_din_pass_2_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_0_6_V_V_full_n_pass_1(fifo_cout_drain_cout_drain_IO_L1_out_0_6_V_V_full_n_pass_1_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_0_6_V_V_full_n_pass_2(fifo_cout_drain_cout_drain_IO_L1_out_0_6_V_V_full_n_pass_2_in),
    .cout_drain_IO_L1_out_wrapper376_U0_fifo_cout_drain_out_V_V_write_pass_1(cout_drain_IO_L1_out_wrapper376_U0_fifo_cout_drain_out_V_V_write_pass_1_in),
    .cout_drain_IO_L1_out_wrapper376_U0_fifo_cout_drain_out_V_V_write_pass_2(cout_drain_IO_L1_out_wrapper376_U0_fifo_cout_drain_out_V_V_write_pass_2_out),
    .PE_wrapper151_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper151_U0_fifo_cout_drain_out_V_din_pass_0_in),
    .PE_wrapper151_U0_fifo_cout_drain_out_V_din_pass_1(PE_wrapper151_U0_fifo_cout_drain_out_V_din_pass_1_out),
    .fifo_cout_drain_PE_0_1_V_full_n_pass_0(fifo_cout_drain_PE_0_1_V_full_n_pass_0_out),
    .fifo_cout_drain_PE_0_1_V_full_n_pass_1(fifo_cout_drain_PE_0_1_V_full_n_pass_1_in),
    .PE_wrapper151_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper151_U0_fifo_cout_drain_out_V_write_pass_0_in),
    .PE_wrapper151_U0_fifo_cout_drain_out_V_write_pass_1(PE_wrapper151_U0_fifo_cout_drain_out_V_write_pass_1_out),
    .cout_drain_IO_L1_out_wrapper392_U0_fifo_cout_drain_out_V_V_din_pass_1(cout_drain_IO_L1_out_wrapper392_U0_fifo_cout_drain_out_V_V_din_pass_1_in),
    .cout_drain_IO_L1_out_wrapper392_U0_fifo_cout_drain_out_V_V_din_pass_2(cout_drain_IO_L1_out_wrapper392_U0_fifo_cout_drain_out_V_V_din_pass_2_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_1_6_V_V_full_n_pass_1(fifo_cout_drain_cout_drain_IO_L1_out_1_6_V_V_full_n_pass_1_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_1_6_V_V_full_n_pass_2(fifo_cout_drain_cout_drain_IO_L1_out_1_6_V_V_full_n_pass_2_in),
    .cout_drain_IO_L1_out_wrapper392_U0_fifo_cout_drain_out_V_V_write_pass_1(cout_drain_IO_L1_out_wrapper392_U0_fifo_cout_drain_out_V_V_write_pass_1_in),
    .cout_drain_IO_L1_out_wrapper392_U0_fifo_cout_drain_out_V_V_write_pass_2(cout_drain_IO_L1_out_wrapper392_U0_fifo_cout_drain_out_V_V_write_pass_2_out),
    .cout_drain_IO_L2_out564_U0_fifo_cout_drain_out_V_V_din_pass_1(cout_drain_IO_L2_out564_U0_fifo_cout_drain_out_V_V_din_pass_1_in),
    .fifo_cout_drain_cout_drain_IO_L2_out_4_V_V_full_n_pass_1(fifo_cout_drain_cout_drain_IO_L2_out_4_V_V_full_n_pass_1_out),
    .cout_drain_IO_L2_out564_U0_fifo_cout_drain_out_V_V_write_pass_1(cout_drain_IO_L2_out564_U0_fifo_cout_drain_out_V_V_write_pass_1_in),
    .PE_wrapper200_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper200_U0_fifo_cout_drain_out_V_din_pass_0_in),
    .fifo_cout_drain_PE_4_2_V_full_n_pass_0(fifo_cout_drain_PE_4_2_V_full_n_pass_0_out),
    .PE_wrapper200_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper200_U0_fifo_cout_drain_out_V_write_pass_0_in),
    .PE_wrapper212_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper212_U0_fifo_cin_out_V_V_din_pass_0_out),
    .fifo_cin_PE_6_2_V_V_full_n_pass_0(fifo_cin_PE_6_2_V_V_full_n_pass_0_in),
    .PE_wrapper212_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper212_U0_fifo_cin_out_V_V_write_pass_0_out),
    .PE_wrapper210_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper210_U0_fifo_w_out_V_V_din_pass_0_in),
    .fifo_w_PE_5_1_V_V_full_n_pass_0(fifo_w_PE_5_1_V_V_full_n_pass_0_out),
    .PE_wrapper210_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper210_U0_fifo_w_out_V_V_write_pass_0_in),
    .PE_wrapper188_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper188_U0_fifo_cout_drain_out_V_din_pass_0_in),
    .fifo_cout_drain_PE_3_2_V_full_n_pass_0(fifo_cout_drain_PE_3_2_V_full_n_pass_0_out),
    .PE_wrapper188_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper188_U0_fifo_cout_drain_out_V_write_pass_0_in),
    .cout_drain_IO_L1_out_wrapper424_U0_fifo_cout_drain_out_V_V_din_pass_1(cout_drain_IO_L1_out_wrapper424_U0_fifo_cout_drain_out_V_V_din_pass_1_in),
    .fifo_cout_drain_cout_drain_IO_L1_out_3_6_V_V_full_n_pass_1(fifo_cout_drain_cout_drain_IO_L1_out_3_6_V_V_full_n_pass_1_out),
    .cout_drain_IO_L1_out_wrapper424_U0_fifo_cout_drain_out_V_V_write_pass_1(cout_drain_IO_L1_out_wrapper424_U0_fifo_cout_drain_out_V_V_write_pass_1_in),
    .PE_wrapper201_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper201_U0_fifo_cin_out_V_V_din_pass_0_in),
    .fifo_cin_PE_5_3_V_V_full_n_pass_0(fifo_cin_PE_5_3_V_V_full_n_pass_0_out),
    .PE_wrapper201_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper201_U0_fifo_cin_out_V_V_write_pass_0_in),
    .cout_drain_IO_L1_out_wrapper398_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper398_U0_fifo_cout_drain_out_V_V_din_pass_0_in),
    .fifo_cout_drain_cout_drain_IO_L1_out_1_0_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_1_0_V_V_full_n_pass_0_out),
    .cout_drain_IO_L1_out_wrapper398_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper398_U0_fifo_cout_drain_out_V_V_write_pass_0_in),
    .PE_wrapper199_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper199_U0_fifo_cin_out_V_V_din_pass_0_in),
    .fifo_cin_PE_5_1_V_V_full_n_pass_0(fifo_cin_PE_5_1_V_V_full_n_pass_0_out),
    .PE_wrapper199_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper199_U0_fifo_cin_out_V_V_write_pass_0_in),
    .PE_wrapper211_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper211_U0_fifo_cin_out_V_V_din_pass_0_out),
    .fifo_cin_PE_6_1_V_V_full_n_pass_0(fifo_cin_PE_6_1_V_V_full_n_pass_0_in),
    .PE_wrapper211_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper211_U0_fifo_cin_out_V_V_write_pass_0_out),
    .PE_wrapper165_U0_fifo_cout_drain_out_V_din_pass_1(PE_wrapper165_U0_fifo_cout_drain_out_V_din_pass_1_in),
    .fifo_cout_drain_PE_1_3_V_full_n_pass_1(fifo_cout_drain_PE_1_3_V_full_n_pass_1_out),
    .PE_wrapper165_U0_fifo_cout_drain_out_V_write_pass_1(PE_wrapper165_U0_fifo_cout_drain_out_V_write_pass_1_in),
    .PE_wrapper211_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper211_U0_fifo_cout_drain_out_V_din_pass_0_out),
    .fifo_cout_drain_PE_5_1_V_full_n_pass_0(fifo_cout_drain_PE_5_1_V_full_n_pass_0_in),
    .PE_wrapper211_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper211_U0_fifo_cout_drain_out_V_write_pass_0_out),
    .PE_wrapper153_U0_fifo_cout_drain_out_V_din_pass_1(PE_wrapper153_U0_fifo_cout_drain_out_V_din_pass_1_in),
    .fifo_cout_drain_PE_0_3_V_full_n_pass_1(fifo_cout_drain_PE_0_3_V_full_n_pass_1_out),
    .PE_wrapper153_U0_fifo_cout_drain_out_V_write_pass_1(PE_wrapper153_U0_fifo_cout_drain_out_V_write_pass_1_in),
    .PE_wrapper201_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper201_U0_fifo_cout_drain_out_V_din_pass_0_in),
    .fifo_cout_drain_PE_4_3_V_full_n_pass_0(fifo_cout_drain_PE_4_3_V_full_n_pass_0_out),
    .PE_wrapper201_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper201_U0_fifo_cout_drain_out_V_write_pass_0_in),
    .cout_drain_IO_L1_out_wrapper382_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper382_U0_fifo_cout_drain_out_V_V_din_pass_0_in),
    .fifo_cout_drain_cout_drain_IO_L1_out_0_0_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_0_0_V_V_full_n_pass_0_out),
    .cout_drain_IO_L1_out_wrapper382_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper382_U0_fifo_cout_drain_out_V_V_write_pass_0_in),
    .PE_wrapper213_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper213_U0_fifo_cin_out_V_V_din_pass_0_out),
    .fifo_cin_PE_6_3_V_V_full_n_pass_0(fifo_cin_PE_6_3_V_V_full_n_pass_0_in),
    .PE_wrapper213_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper213_U0_fifo_cin_out_V_V_write_pass_0_out),
    .PE_wrapper177_U0_fifo_cout_drain_out_V_din_pass_1(PE_wrapper177_U0_fifo_cout_drain_out_V_din_pass_1_in),
    .fifo_cout_drain_PE_2_3_V_full_n_pass_1(fifo_cout_drain_PE_2_3_V_full_n_pass_1_out),
    .PE_wrapper177_U0_fifo_cout_drain_out_V_write_pass_1(PE_wrapper177_U0_fifo_cout_drain_out_V_write_pass_1_in),
    .PE_wrapper164_U0_fifo_cout_drain_out_V_din_pass_1(PE_wrapper164_U0_fifo_cout_drain_out_V_din_pass_1_in),
    .fifo_cout_drain_PE_1_2_V_full_n_pass_1(fifo_cout_drain_PE_1_2_V_full_n_pass_1_out),
    .PE_wrapper164_U0_fifo_cout_drain_out_V_write_pass_1(PE_wrapper164_U0_fifo_cout_drain_out_V_write_pass_1_in),
    .PE_wrapper189_U0_fifo_cout_drain_out_V_din_pass_1(PE_wrapper189_U0_fifo_cout_drain_out_V_din_pass_1_in),
    .fifo_cout_drain_PE_3_3_V_full_n_pass_1(fifo_cout_drain_PE_3_3_V_full_n_pass_1_out),
    .PE_wrapper189_U0_fifo_cout_drain_out_V_write_pass_1(PE_wrapper189_U0_fifo_cout_drain_out_V_write_pass_1_in),
    .cin_IO_L2_in124_U0_fifo_cin_out_V_V_din_pass_0(cin_IO_L2_in124_U0_fifo_cin_out_V_V_din_pass_0_in),
    .fifo_cin_cin_IO_L2_in_1_V_V_full_n_pass_0(fifo_cin_cin_IO_L2_in_1_V_V_full_n_pass_0_out),
    .cin_IO_L2_in124_U0_fifo_cin_out_V_V_write_pass_0(cin_IO_L2_in124_U0_fifo_cin_out_V_V_write_pass_0_in),
    .PE_wrapper152_U0_fifo_cout_drain_out_V_din_pass_1(PE_wrapper152_U0_fifo_cout_drain_out_V_din_pass_1_in),
    .fifo_cout_drain_PE_0_2_V_full_n_pass_1(fifo_cout_drain_PE_0_2_V_full_n_pass_1_out),
    .PE_wrapper152_U0_fifo_cout_drain_out_V_write_pass_1(PE_wrapper152_U0_fifo_cout_drain_out_V_write_pass_1_in),
    .cin_IO_L2_in125_U0_fifo_cin_out_V_V_din_pass_0(cin_IO_L2_in125_U0_fifo_cin_out_V_V_din_pass_0_out),
    .fifo_cin_cin_IO_L2_in_2_V_V_full_n_pass_0(fifo_cin_cin_IO_L2_in_2_V_V_full_n_pass_0_in),
    .cin_IO_L2_in125_U0_fifo_cin_out_V_V_write_pass_0(cin_IO_L2_in125_U0_fifo_cin_out_V_V_write_pass_0_out),
    .PE_wrapper200_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper200_U0_fifo_cin_out_V_V_din_pass_0_in),
    .fifo_cin_PE_5_2_V_V_full_n_pass_0(fifo_cin_PE_5_2_V_V_full_n_pass_0_out),
    .PE_wrapper200_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper200_U0_fifo_cin_out_V_V_write_pass_0_in),
    .cin_IO_L2_in125_U0_fifo_cin_local_out_V_V_din_pass_0(cin_IO_L2_in125_U0_fifo_cin_local_out_V_V_din_pass_0_out),
    .fifo_cin_PE_0_1_V_V_full_n_pass_0(fifo_cin_PE_0_1_V_V_full_n_pass_0_in),
    .cin_IO_L2_in125_U0_fifo_cin_local_out_V_V_write_pass_0(cin_IO_L2_in125_U0_fifo_cin_local_out_V_V_write_pass_0_out),
    .cout_drain_IO_L1_out_wrapper408_U0_fifo_cout_drain_out_V_V_din_pass_1(cout_drain_IO_L1_out_wrapper408_U0_fifo_cout_drain_out_V_V_din_pass_1_in),
    .fifo_cout_drain_cout_drain_IO_L1_out_2_6_V_V_full_n_pass_1(fifo_cout_drain_cout_drain_IO_L1_out_2_6_V_V_full_n_pass_1_out),
    .cout_drain_IO_L1_out_wrapper408_U0_fifo_cout_drain_out_V_V_write_pass_1(cout_drain_IO_L1_out_wrapper408_U0_fifo_cout_drain_out_V_V_write_pass_1_in),
    .PE_wrapper213_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper213_U0_fifo_w_out_V_V_din_pass_0_out),
    .fifo_w_PE_5_4_V_V_full_n_pass_0(fifo_w_PE_5_4_V_V_full_n_pass_0_in),
    .PE_wrapper213_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper213_U0_fifo_w_out_V_V_write_pass_0_out),
    .cout_drain_IO_L2_out568_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L2_out568_U0_fifo_cout_drain_out_V_V_din_pass_0_out),
    .fifo_cout_drain_cout_drain_IO_L2_out_0_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L2_out_0_V_V_full_n_pass_0_in),
    .cout_drain_IO_L2_out568_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L2_out568_U0_fifo_cout_drain_out_V_V_write_pass_0_out),
    .PE_wrapper176_U0_fifo_cout_drain_out_V_din_pass_1(PE_wrapper176_U0_fifo_cout_drain_out_V_din_pass_1_in),
    .fifo_cout_drain_PE_2_2_V_full_n_pass_1(fifo_cout_drain_PE_2_2_V_full_n_pass_1_out),
    .PE_wrapper176_U0_fifo_cout_drain_out_V_write_pass_1(PE_wrapper176_U0_fifo_cout_drain_out_V_write_pass_1_in),
    .ap_clk(ap_clk),
    .ap_start_Boundary_X6Y0_To_X6Y2(ap_start_Boundary_X6Y0_To_X6Y2_in),
    .ap_rst_n_Boundary_X6Y0_To_X6Y2(ap_rst_n_Boundary_X6Y0_To_X6Y2_in),
    .ap_done_Boundary_X6Y0_To_X6Y2(ap_done_Boundary_X6Y0_To_X6Y2_out),
    .ap_start_Boundary_X6Y2_To_X8Y2(ap_start_Boundary_X6Y2_To_X8Y2_out),
    .ap_rst_n_Boundary_X6Y2_To_X8Y2(ap_rst_n_Boundary_X6Y2_To_X8Y2_out),
    .ap_done_Boundary_X6Y2_To_X8Y2(ap_done_Boundary_X6Y2_To_X8Y2_in)
  );


  (* keep_hierarchy = "yes" *) CR_X6Y2_To_CR_X7Y3_ctrl CR_X6Y2_To_CR_X7Y3_ctrl_U0 (
    .cout_drain_IO_L2_out564_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L2_out564_U0_fifo_cout_drain_out_V_V_din_pass_0_in),
    .cout_drain_IO_L2_out564_U0_fifo_cout_drain_out_V_V_din_pass_1(cout_drain_IO_L2_out564_U0_fifo_cout_drain_out_V_V_din_pass_1_out),
    .fifo_cout_drain_cout_drain_IO_L2_out_4_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L2_out_4_V_V_full_n_pass_0_out),
    .fifo_cout_drain_cout_drain_IO_L2_out_4_V_V_full_n_pass_1(fifo_cout_drain_cout_drain_IO_L2_out_4_V_V_full_n_pass_1_in),
    .cout_drain_IO_L2_out564_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L2_out564_U0_fifo_cout_drain_out_V_V_write_pass_0_in),
    .cout_drain_IO_L2_out564_U0_fifo_cout_drain_out_V_V_write_pass_1(cout_drain_IO_L2_out564_U0_fifo_cout_drain_out_V_V_write_pass_1_out),
    .PE_wrapper165_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper165_U0_fifo_cout_drain_out_V_din_pass_0_in),
    .PE_wrapper165_U0_fifo_cout_drain_out_V_din_pass_1(PE_wrapper165_U0_fifo_cout_drain_out_V_din_pass_1_out),
    .fifo_cout_drain_PE_1_3_V_full_n_pass_0(fifo_cout_drain_PE_1_3_V_full_n_pass_0_out),
    .fifo_cout_drain_PE_1_3_V_full_n_pass_1(fifo_cout_drain_PE_1_3_V_full_n_pass_1_in),
    .PE_wrapper165_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper165_U0_fifo_cout_drain_out_V_write_pass_0_in),
    .PE_wrapper165_U0_fifo_cout_drain_out_V_write_pass_1(PE_wrapper165_U0_fifo_cout_drain_out_V_write_pass_1_out),
    .PE_wrapper153_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper153_U0_fifo_cout_drain_out_V_din_pass_0_in),
    .PE_wrapper153_U0_fifo_cout_drain_out_V_din_pass_1(PE_wrapper153_U0_fifo_cout_drain_out_V_din_pass_1_out),
    .fifo_cout_drain_PE_0_3_V_full_n_pass_0(fifo_cout_drain_PE_0_3_V_full_n_pass_0_out),
    .fifo_cout_drain_PE_0_3_V_full_n_pass_1(fifo_cout_drain_PE_0_3_V_full_n_pass_1_in),
    .PE_wrapper153_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper153_U0_fifo_cout_drain_out_V_write_pass_0_in),
    .PE_wrapper153_U0_fifo_cout_drain_out_V_write_pass_1(PE_wrapper153_U0_fifo_cout_drain_out_V_write_pass_1_out),
    .PE_wrapper177_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper177_U0_fifo_cout_drain_out_V_din_pass_0_in),
    .PE_wrapper177_U0_fifo_cout_drain_out_V_din_pass_1(PE_wrapper177_U0_fifo_cout_drain_out_V_din_pass_1_out),
    .fifo_cout_drain_PE_2_3_V_full_n_pass_0(fifo_cout_drain_PE_2_3_V_full_n_pass_0_out),
    .fifo_cout_drain_PE_2_3_V_full_n_pass_1(fifo_cout_drain_PE_2_3_V_full_n_pass_1_in),
    .PE_wrapper177_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper177_U0_fifo_cout_drain_out_V_write_pass_0_in),
    .PE_wrapper177_U0_fifo_cout_drain_out_V_write_pass_1(PE_wrapper177_U0_fifo_cout_drain_out_V_write_pass_1_out),
    .PE_wrapper164_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper164_U0_fifo_cout_drain_out_V_din_pass_0_in),
    .PE_wrapper164_U0_fifo_cout_drain_out_V_din_pass_1(PE_wrapper164_U0_fifo_cout_drain_out_V_din_pass_1_out),
    .fifo_cout_drain_PE_1_2_V_full_n_pass_0(fifo_cout_drain_PE_1_2_V_full_n_pass_0_out),
    .fifo_cout_drain_PE_1_2_V_full_n_pass_1(fifo_cout_drain_PE_1_2_V_full_n_pass_1_in),
    .PE_wrapper164_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper164_U0_fifo_cout_drain_out_V_write_pass_0_in),
    .PE_wrapper164_U0_fifo_cout_drain_out_V_write_pass_1(PE_wrapper164_U0_fifo_cout_drain_out_V_write_pass_1_out),
    .PE_wrapper189_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper189_U0_fifo_cout_drain_out_V_din_pass_0_in),
    .PE_wrapper189_U0_fifo_cout_drain_out_V_din_pass_1(PE_wrapper189_U0_fifo_cout_drain_out_V_din_pass_1_out),
    .fifo_cout_drain_PE_3_3_V_full_n_pass_0(fifo_cout_drain_PE_3_3_V_full_n_pass_0_out),
    .fifo_cout_drain_PE_3_3_V_full_n_pass_1(fifo_cout_drain_PE_3_3_V_full_n_pass_1_in),
    .PE_wrapper189_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper189_U0_fifo_cout_drain_out_V_write_pass_0_in),
    .PE_wrapper189_U0_fifo_cout_drain_out_V_write_pass_1(PE_wrapper189_U0_fifo_cout_drain_out_V_write_pass_1_out),
    .PE_wrapper152_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper152_U0_fifo_cout_drain_out_V_din_pass_0_in),
    .PE_wrapper152_U0_fifo_cout_drain_out_V_din_pass_1(PE_wrapper152_U0_fifo_cout_drain_out_V_din_pass_1_out),
    .fifo_cout_drain_PE_0_2_V_full_n_pass_0(fifo_cout_drain_PE_0_2_V_full_n_pass_0_out),
    .fifo_cout_drain_PE_0_2_V_full_n_pass_1(fifo_cout_drain_PE_0_2_V_full_n_pass_1_in),
    .PE_wrapper152_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper152_U0_fifo_cout_drain_out_V_write_pass_0_in),
    .PE_wrapper152_U0_fifo_cout_drain_out_V_write_pass_1(PE_wrapper152_U0_fifo_cout_drain_out_V_write_pass_1_out),
    .PE_wrapper176_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper176_U0_fifo_cout_drain_out_V_din_pass_0_in),
    .PE_wrapper176_U0_fifo_cout_drain_out_V_din_pass_1(PE_wrapper176_U0_fifo_cout_drain_out_V_din_pass_1_out),
    .fifo_cout_drain_PE_2_2_V_full_n_pass_0(fifo_cout_drain_PE_2_2_V_full_n_pass_0_out),
    .fifo_cout_drain_PE_2_2_V_full_n_pass_1(fifo_cout_drain_PE_2_2_V_full_n_pass_1_in),
    .PE_wrapper176_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper176_U0_fifo_cout_drain_out_V_write_pass_0_in),
    .PE_wrapper176_U0_fifo_cout_drain_out_V_write_pass_1(PE_wrapper176_U0_fifo_cout_drain_out_V_write_pass_1_out),
    .PE_wrapper165_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper165_U0_fifo_w_out_V_V_din_pass_0_in),
    .PE_wrapper165_U0_fifo_w_out_V_V_din_pass_1(PE_wrapper165_U0_fifo_w_out_V_V_din_pass_1_out),
    .fifo_w_PE_1_4_V_V_full_n_pass_0(fifo_w_PE_1_4_V_V_full_n_pass_0_out),
    .fifo_w_PE_1_4_V_V_full_n_pass_1(fifo_w_PE_1_4_V_V_full_n_pass_1_in),
    .PE_wrapper165_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper165_U0_fifo_w_out_V_V_write_pass_0_in),
    .PE_wrapper165_U0_fifo_w_out_V_V_write_pass_1(PE_wrapper165_U0_fifo_w_out_V_V_write_pass_1_out),
    .cin_IO_L2_in127_U0_fifo_cin_out_V_V_din_pass_0(cin_IO_L2_in127_U0_fifo_cin_out_V_V_din_pass_0_in),
    .cin_IO_L2_in127_U0_fifo_cin_out_V_V_din_pass_1(cin_IO_L2_in127_U0_fifo_cin_out_V_V_din_pass_1_out),
    .fifo_cin_cin_IO_L2_in_4_V_V_full_n_pass_0(fifo_cin_cin_IO_L2_in_4_V_V_full_n_pass_0_out),
    .fifo_cin_cin_IO_L2_in_4_V_V_full_n_pass_1(fifo_cin_cin_IO_L2_in_4_V_V_full_n_pass_1_in),
    .cin_IO_L2_in127_U0_fifo_cin_out_V_V_write_pass_0(cin_IO_L2_in127_U0_fifo_cin_out_V_V_write_pass_0_in),
    .cin_IO_L2_in127_U0_fifo_cin_out_V_V_write_pass_1(cin_IO_L2_in127_U0_fifo_cin_out_V_V_write_pass_1_out),
    .PE_wrapper177_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper177_U0_fifo_w_out_V_V_din_pass_0_in),
    .PE_wrapper177_U0_fifo_w_out_V_V_din_pass_1(PE_wrapper177_U0_fifo_w_out_V_V_din_pass_1_out),
    .fifo_w_PE_2_4_V_V_full_n_pass_0(fifo_w_PE_2_4_V_V_full_n_pass_0_out),
    .fifo_w_PE_2_4_V_V_full_n_pass_1(fifo_w_PE_2_4_V_V_full_n_pass_1_in),
    .PE_wrapper177_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper177_U0_fifo_w_out_V_V_write_pass_0_in),
    .PE_wrapper177_U0_fifo_w_out_V_V_write_pass_1(PE_wrapper177_U0_fifo_w_out_V_V_write_pass_1_out),
    .PE_wrapper153_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper153_U0_fifo_w_out_V_V_din_pass_0_in),
    .PE_wrapper153_U0_fifo_w_out_V_V_din_pass_1(PE_wrapper153_U0_fifo_w_out_V_V_din_pass_1_out),
    .fifo_w_PE_0_4_V_V_full_n_pass_0(fifo_w_PE_0_4_V_V_full_n_pass_0_out),
    .fifo_w_PE_0_4_V_V_full_n_pass_1(fifo_w_PE_0_4_V_V_full_n_pass_1_in),
    .PE_wrapper153_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper153_U0_fifo_w_out_V_V_write_pass_0_in),
    .PE_wrapper153_U0_fifo_w_out_V_V_write_pass_1(PE_wrapper153_U0_fifo_w_out_V_V_write_pass_1_out),
    .PE_wrapper189_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper189_U0_fifo_w_out_V_V_din_pass_0_in),
    .PE_wrapper189_U0_fifo_w_out_V_V_din_pass_1(PE_wrapper189_U0_fifo_w_out_V_V_din_pass_1_out),
    .fifo_w_PE_3_4_V_V_full_n_pass_0(fifo_w_PE_3_4_V_V_full_n_pass_0_out),
    .fifo_w_PE_3_4_V_V_full_n_pass_1(fifo_w_PE_3_4_V_V_full_n_pass_1_in),
    .PE_wrapper189_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper189_U0_fifo_w_out_V_V_write_pass_0_in),
    .PE_wrapper189_U0_fifo_w_out_V_V_write_pass_1(PE_wrapper189_U0_fifo_w_out_V_V_write_pass_1_out),
    .cout_drain_IO_L2_out568_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L2_out568_U0_fifo_cout_drain_out_V_V_din_pass_0_in),
    .cout_drain_IO_L2_out568_U0_fifo_cout_drain_out_V_V_din_pass_1(cout_drain_IO_L2_out568_U0_fifo_cout_drain_out_V_V_din_pass_1_out),
    .fifo_cout_drain_cout_drain_IO_L2_out_0_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L2_out_0_V_V_full_n_pass_0_out),
    .fifo_cout_drain_cout_drain_IO_L2_out_0_V_V_full_n_pass_1(fifo_cout_drain_cout_drain_IO_L2_out_0_V_V_full_n_pass_1_in),
    .cout_drain_IO_L2_out568_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L2_out568_U0_fifo_cout_drain_out_V_V_write_pass_0_in),
    .cout_drain_IO_L2_out568_U0_fifo_cout_drain_out_V_V_write_pass_1(cout_drain_IO_L2_out568_U0_fifo_cout_drain_out_V_V_write_pass_1_out),
    .w_IO_L2_in140_U0_fifo_w_out_V_V_din_pass_0(w_IO_L2_in140_U0_fifo_w_out_V_V_din_pass_0_out),
    .fifo_w_w_IO_L2_in_6_V_V_full_n_pass_0(fifo_w_w_IO_L2_in_6_V_V_full_n_pass_0_in),
    .w_IO_L2_in140_U0_fifo_w_out_V_V_write_pass_0(w_IO_L2_in140_U0_fifo_w_out_V_V_write_pass_0_out),
    .PE_wrapper187_U0_fifo_w_out_V_V_din_pass_1(PE_wrapper187_U0_fifo_w_out_V_V_din_pass_1_in),
    .fifo_w_PE_3_2_V_V_full_n_pass_1(fifo_w_PE_3_2_V_V_full_n_pass_1_out),
    .PE_wrapper187_U0_fifo_w_out_V_V_write_pass_1(PE_wrapper187_U0_fifo_w_out_V_V_write_pass_1_in),
    .PE_wrapper188_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper188_U0_fifo_w_out_V_V_din_pass_0_out),
    .fifo_w_PE_3_3_V_V_full_n_pass_0(fifo_w_PE_3_3_V_V_full_n_pass_0_in),
    .PE_wrapper188_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper188_U0_fifo_w_out_V_V_write_pass_0_out),
    .PE_wrapper200_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper200_U0_fifo_cout_drain_out_V_din_pass_0_out),
    .fifo_cout_drain_PE_4_2_V_full_n_pass_0(fifo_cout_drain_PE_4_2_V_full_n_pass_0_in),
    .PE_wrapper200_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper200_U0_fifo_cout_drain_out_V_write_pass_0_out),
    .PE_wrapper188_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper188_U0_fifo_cout_drain_out_V_din_pass_0_out),
    .fifo_cout_drain_PE_3_2_V_full_n_pass_0(fifo_cout_drain_PE_3_2_V_full_n_pass_0_in),
    .PE_wrapper188_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper188_U0_fifo_cout_drain_out_V_write_pass_0_out),
    .PE_wrapper210_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper210_U0_fifo_w_out_V_V_din_pass_0_out),
    .fifo_w_PE_5_1_V_V_full_n_pass_0(fifo_w_PE_5_1_V_V_full_n_pass_0_in),
    .PE_wrapper210_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper210_U0_fifo_w_out_V_V_write_pass_0_out),
    .PE_wrapper201_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper201_U0_fifo_cin_out_V_V_din_pass_0_out),
    .fifo_cin_PE_5_3_V_V_full_n_pass_0(fifo_cin_PE_5_3_V_V_full_n_pass_0_in),
    .PE_wrapper201_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper201_U0_fifo_cin_out_V_V_write_pass_0_out),
    .cout_drain_IO_L1_out_wrapper398_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper398_U0_fifo_cout_drain_out_V_V_din_pass_0_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_1_0_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_1_0_V_V_full_n_pass_0_in),
    .cout_drain_IO_L1_out_wrapper398_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper398_U0_fifo_cout_drain_out_V_V_write_pass_0_out),
    .PE_wrapper199_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper199_U0_fifo_cin_out_V_V_din_pass_0_out),
    .fifo_cin_PE_5_1_V_V_full_n_pass_0(fifo_cin_PE_5_1_V_V_full_n_pass_0_in),
    .PE_wrapper199_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper199_U0_fifo_cin_out_V_V_write_pass_0_out),
    .PE_wrapper163_U0_fifo_cout_drain_out_V_din_pass_1(PE_wrapper163_U0_fifo_cout_drain_out_V_din_pass_1_in),
    .fifo_cout_drain_PE_1_1_V_full_n_pass_1(fifo_cout_drain_PE_1_1_V_full_n_pass_1_out),
    .PE_wrapper163_U0_fifo_cout_drain_out_V_write_pass_1(PE_wrapper163_U0_fifo_cout_drain_out_V_write_pass_1_in),
    .PE_wrapper211_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper211_U0_fifo_cout_drain_out_V_din_pass_0_in),
    .fifo_cout_drain_PE_5_1_V_full_n_pass_0(fifo_cout_drain_PE_5_1_V_full_n_pass_0_out),
    .PE_wrapper211_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper211_U0_fifo_cout_drain_out_V_write_pass_0_in),
    .cout_drain_IO_L1_out_wrapper378_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper378_U0_fifo_cout_drain_out_V_V_din_pass_0_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_0_4_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_0_4_V_V_full_n_pass_0_in),
    .cout_drain_IO_L1_out_wrapper378_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper378_U0_fifo_cout_drain_out_V_V_write_pass_0_out),
    .PE_wrapper175_U0_fifo_cout_drain_out_V_din_pass_1(PE_wrapper175_U0_fifo_cout_drain_out_V_din_pass_1_in),
    .fifo_cout_drain_PE_2_1_V_full_n_pass_1(fifo_cout_drain_PE_2_1_V_full_n_pass_1_out),
    .PE_wrapper175_U0_fifo_cout_drain_out_V_write_pass_1(PE_wrapper175_U0_fifo_cout_drain_out_V_write_pass_1_in),
    .PE_wrapper201_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper201_U0_fifo_cout_drain_out_V_din_pass_0_out),
    .fifo_cout_drain_PE_4_3_V_full_n_pass_0(fifo_cout_drain_PE_4_3_V_full_n_pass_0_in),
    .PE_wrapper201_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper201_U0_fifo_cout_drain_out_V_write_pass_0_out),
    .PE_wrapper187_U0_fifo_cin_out_V_V_din_pass_1(PE_wrapper187_U0_fifo_cin_out_V_V_din_pass_1_in),
    .fifo_cin_PE_4_1_V_V_full_n_pass_1(fifo_cin_PE_4_1_V_V_full_n_pass_1_out),
    .PE_wrapper187_U0_fifo_cin_out_V_V_write_pass_1(PE_wrapper187_U0_fifo_cin_out_V_V_write_pass_1_in),
    .PE_wrapper186_U0_fifo_cin_out_V_V_din_pass_1(PE_wrapper186_U0_fifo_cin_out_V_V_din_pass_1_in),
    .fifo_cin_PE_4_0_V_V_full_n_pass_1(fifo_cin_PE_4_0_V_V_full_n_pass_1_out),
    .PE_wrapper186_U0_fifo_cin_out_V_V_write_pass_1(PE_wrapper186_U0_fifo_cin_out_V_V_write_pass_1_in),
    .PE_wrapper201_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper201_U0_fifo_w_out_V_V_din_pass_0_out),
    .fifo_w_PE_4_4_V_V_full_n_pass_0(fifo_w_PE_4_4_V_V_full_n_pass_0_in),
    .PE_wrapper201_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper201_U0_fifo_w_out_V_V_write_pass_0_out),
    .PE_wrapper187_U0_fifo_cout_drain_out_V_din_pass_1(PE_wrapper187_U0_fifo_cout_drain_out_V_din_pass_1_in),
    .fifo_cout_drain_PE_3_1_V_full_n_pass_1(fifo_cout_drain_PE_3_1_V_full_n_pass_1_out),
    .PE_wrapper187_U0_fifo_cout_drain_out_V_write_pass_1(PE_wrapper187_U0_fifo_cout_drain_out_V_write_pass_1_in),
    .w_IO_L2_in137_U0_fifo_w_out_V_V_din_pass_1(w_IO_L2_in137_U0_fifo_w_out_V_V_din_pass_1_in),
    .fifo_w_w_IO_L2_in_3_V_V_full_n_pass_1(fifo_w_w_IO_L2_in_3_V_V_full_n_pass_1_out),
    .w_IO_L2_in137_U0_fifo_w_out_V_V_write_pass_1(w_IO_L2_in137_U0_fifo_w_out_V_V_write_pass_1_in),
    .cout_drain_IO_L1_out_wrapper376_U0_fifo_cout_drain_out_V_V_din_pass_2(cout_drain_IO_L1_out_wrapper376_U0_fifo_cout_drain_out_V_V_din_pass_2_in),
    .fifo_cout_drain_cout_drain_IO_L1_out_0_6_V_V_full_n_pass_2(fifo_cout_drain_cout_drain_IO_L1_out_0_6_V_V_full_n_pass_2_out),
    .cout_drain_IO_L1_out_wrapper376_U0_fifo_cout_drain_out_V_V_write_pass_2(cout_drain_IO_L1_out_wrapper376_U0_fifo_cout_drain_out_V_V_write_pass_2_in),
    .PE_wrapper151_U0_fifo_cout_drain_out_V_din_pass_1(PE_wrapper151_U0_fifo_cout_drain_out_V_din_pass_1_in),
    .fifo_cout_drain_PE_0_1_V_full_n_pass_1(fifo_cout_drain_PE_0_1_V_full_n_pass_1_out),
    .PE_wrapper151_U0_fifo_cout_drain_out_V_write_pass_1(PE_wrapper151_U0_fifo_cout_drain_out_V_write_pass_1_in),
    .w_IO_L2_in138_U0_fifo_w_local_out_V_V_din_pass_0(w_IO_L2_in138_U0_fifo_w_local_out_V_V_din_pass_0_out),
    .fifo_w_PE_3_0_V_V_full_n_pass_0(fifo_w_PE_3_0_V_V_full_n_pass_0_in),
    .w_IO_L2_in138_U0_fifo_w_local_out_V_V_write_pass_0(w_IO_L2_in138_U0_fifo_w_local_out_V_V_write_pass_0_out),
    .PE_wrapper200_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper200_U0_fifo_cin_out_V_V_din_pass_0_out),
    .fifo_cin_PE_5_2_V_V_full_n_pass_0(fifo_cin_PE_5_2_V_V_full_n_pass_0_in),
    .PE_wrapper200_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper200_U0_fifo_cin_out_V_V_write_pass_0_out),
    .PE_wrapper189_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper189_U0_fifo_cin_out_V_V_din_pass_0_in),
    .fifo_cin_PE_4_3_V_V_full_n_pass_0(fifo_cin_PE_4_3_V_V_full_n_pass_0_out),
    .PE_wrapper189_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper189_U0_fifo_cin_out_V_V_write_pass_0_in),
    .PE_wrapper176_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper176_U0_fifo_cin_out_V_V_din_pass_0_in),
    .fifo_cin_PE_3_2_V_V_full_n_pass_0(fifo_cin_PE_3_2_V_V_full_n_pass_0_out),
    .PE_wrapper176_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper176_U0_fifo_cin_out_V_V_write_pass_0_in),
    .PE_wrapper210_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper210_U0_fifo_cin_out_V_V_din_pass_0_out),
    .fifo_cin_PE_6_0_V_V_full_n_pass_0(fifo_cin_PE_6_0_V_V_full_n_pass_0_in),
    .PE_wrapper210_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper210_U0_fifo_cin_out_V_V_write_pass_0_out),
    .cout_drain_IO_L1_out_wrapper392_U0_fifo_cout_drain_out_V_V_din_pass_2(cout_drain_IO_L1_out_wrapper392_U0_fifo_cout_drain_out_V_V_din_pass_2_in),
    .fifo_cout_drain_cout_drain_IO_L1_out_1_6_V_V_full_n_pass_2(fifo_cout_drain_cout_drain_IO_L1_out_1_6_V_V_full_n_pass_2_out),
    .cout_drain_IO_L1_out_wrapper392_U0_fifo_cout_drain_out_V_V_write_pass_2(cout_drain_IO_L1_out_wrapper392_U0_fifo_cout_drain_out_V_V_write_pass_2_in),
    .ap_clk(ap_clk),
    .ap_start_Boundary_X6Y2_To_X8Y2(ap_start_Boundary_X6Y2_To_X8Y2_in),
    .ap_rst_n_Boundary_X6Y2_To_X8Y2(ap_rst_n_Boundary_X6Y2_To_X8Y2_in),
    .ap_done_Boundary_X6Y2_To_X8Y2(ap_done_Boundary_X6Y2_To_X8Y2_out),
    .ap_start_Boundary_X6Y4_To_X8Y4(ap_start_Boundary_X6Y4_To_X8Y4_out),
    .ap_rst_n_Boundary_X6Y4_To_X8Y4(ap_rst_n_Boundary_X6Y4_To_X8Y4_out),
    .ap_done_Boundary_X6Y4_To_X8Y4(ap_done_Boundary_X6Y4_To_X8Y4_in)
  );


  (* keep_hierarchy = "yes" *) CR_X4Y6_To_CR_X5Y7_ctrl CR_X4Y6_To_CR_X5Y7_ctrl_U0 (
    .PE_wrapper214_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper214_U0_fifo_w_out_V_V_din_pass_0_in),
    .PE_wrapper214_U0_fifo_w_out_V_V_din_pass_1(PE_wrapper214_U0_fifo_w_out_V_V_din_pass_1_out),
    .fifo_w_PE_5_5_V_V_full_n_pass_0(fifo_w_PE_5_5_V_V_full_n_pass_0_out),
    .fifo_w_PE_5_5_V_V_full_n_pass_1(fifo_w_PE_5_5_V_V_full_n_pass_1_in),
    .PE_wrapper214_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper214_U0_fifo_w_out_V_V_write_pass_0_in),
    .PE_wrapper214_U0_fifo_w_out_V_V_write_pass_1(PE_wrapper214_U0_fifo_w_out_V_V_write_pass_1_out),
    .PE_wrapper202_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper202_U0_fifo_w_out_V_V_din_pass_0_in),
    .PE_wrapper202_U0_fifo_w_out_V_V_din_pass_1(PE_wrapper202_U0_fifo_w_out_V_V_din_pass_1_out),
    .fifo_w_PE_4_5_V_V_full_n_pass_0(fifo_w_PE_4_5_V_V_full_n_pass_0_out),
    .fifo_w_PE_4_5_V_V_full_n_pass_1(fifo_w_PE_4_5_V_V_full_n_pass_1_in),
    .PE_wrapper202_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper202_U0_fifo_w_out_V_V_write_pass_0_in),
    .PE_wrapper202_U0_fifo_w_out_V_V_write_pass_1(PE_wrapper202_U0_fifo_w_out_V_V_write_pass_1_out),
    .kernel0_entry12_U0_cout_V_out_din_pass_2(kernel0_entry12_U0_cout_V_out_din_pass_2_in),
    .kernel0_entry12_U0_cout_V_out_din_pass_3(kernel0_entry12_U0_cout_V_out_din_pass_3_out),
    .cout_V_c_full_n_pass_2(cout_V_c_full_n_pass_2_out),
    .cout_V_c_full_n_pass_3(cout_V_c_full_n_pass_3_in),
    .kernel0_entry12_U0_cout_V_out_write_pass_2(kernel0_entry12_U0_cout_V_out_write_pass_2_in),
    .kernel0_entry12_U0_cout_V_out_write_pass_3(kernel0_entry12_U0_cout_V_out_write_pass_3_out),
    .PE_wrapper243_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper243_U0_fifo_w_out_V_V_din_pass_0_in),
    .PE_wrapper243_U0_fifo_w_out_V_V_din_pass_1(PE_wrapper243_U0_fifo_w_out_V_V_din_pass_1_out),
    .fifo_w_PE_7_10_V_V_full_n_pass_0(fifo_w_PE_7_10_V_V_full_n_pass_0_out),
    .fifo_w_PE_7_10_V_V_full_n_pass_1(fifo_w_PE_7_10_V_V_full_n_pass_1_in),
    .PE_wrapper243_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper243_U0_fifo_w_out_V_V_write_pass_0_in),
    .PE_wrapper243_U0_fifo_w_out_V_V_write_pass_1(PE_wrapper243_U0_fifo_w_out_V_V_write_pass_1_out),
    .PE_wrapper243_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper243_U0_fifo_cout_drain_out_V_din_pass_0_in),
    .PE_wrapper243_U0_fifo_cout_drain_out_V_din_pass_1(PE_wrapper243_U0_fifo_cout_drain_out_V_din_pass_1_out),
    .fifo_cout_drain_PE_7_9_V_full_n_pass_0(fifo_cout_drain_PE_7_9_V_full_n_pass_0_out),
    .fifo_cout_drain_PE_7_9_V_full_n_pass_1(fifo_cout_drain_PE_7_9_V_full_n_pass_1_in),
    .PE_wrapper243_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper243_U0_fifo_cout_drain_out_V_write_pass_0_in),
    .PE_wrapper243_U0_fifo_cout_drain_out_V_write_pass_1(PE_wrapper243_U0_fifo_cout_drain_out_V_write_pass_1_out),
    .PE_wrapper243_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper243_U0_fifo_cin_out_V_V_din_pass_0_in),
    .PE_wrapper243_U0_fifo_cin_out_V_V_din_pass_1(PE_wrapper243_U0_fifo_cin_out_V_V_din_pass_1_out),
    .fifo_cin_PE_8_9_V_V_full_n_pass_0(fifo_cin_PE_8_9_V_V_full_n_pass_0_out),
    .fifo_cin_PE_8_9_V_V_full_n_pass_1(fifo_cin_PE_8_9_V_V_full_n_pass_1_in),
    .PE_wrapper243_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper243_U0_fifo_cin_out_V_V_write_pass_0_in),
    .PE_wrapper243_U0_fifo_cin_out_V_V_write_pass_1(PE_wrapper243_U0_fifo_cin_out_V_V_write_pass_1_out),
    .PE_wrapper191_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper191_U0_fifo_cin_out_V_V_din_pass_0_out),
    .fifo_cin_PE_4_5_V_V_full_n_pass_0(fifo_cin_PE_4_5_V_V_full_n_pass_0_in),
    .PE_wrapper191_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper191_U0_fifo_cin_out_V_V_write_pass_0_out),
    .PE_wrapper191_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper191_U0_fifo_cout_drain_out_V_din_pass_0_out),
    .fifo_cout_drain_PE_3_5_V_full_n_pass_0(fifo_cout_drain_PE_3_5_V_full_n_pass_0_in),
    .PE_wrapper191_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper191_U0_fifo_cout_drain_out_V_write_pass_0_out),
    .PE_wrapper192_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper192_U0_fifo_cin_out_V_V_din_pass_0_out),
    .fifo_cin_PE_4_6_V_V_full_n_pass_0(fifo_cin_PE_4_6_V_V_full_n_pass_0_in),
    .PE_wrapper192_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper192_U0_fifo_cin_out_V_V_write_pass_0_out),
    .PE_wrapper192_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper192_U0_fifo_cout_drain_out_V_din_pass_0_out),
    .fifo_cout_drain_PE_3_6_V_full_n_pass_0(fifo_cout_drain_PE_3_6_V_full_n_pass_0_in),
    .PE_wrapper192_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper192_U0_fifo_cout_drain_out_V_write_pass_0_out),
    .PE_wrapper192_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper192_U0_fifo_w_out_V_V_din_pass_0_out),
    .fifo_w_PE_3_7_V_V_full_n_pass_0(fifo_w_PE_3_7_V_V_full_n_pass_0_in),
    .PE_wrapper192_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper192_U0_fifo_w_out_V_V_write_pass_0_out),
    .PE_wrapper190_U0_fifo_w_out_V_V_din_pass_1(PE_wrapper190_U0_fifo_w_out_V_V_din_pass_1_in),
    .fifo_w_PE_3_5_V_V_full_n_pass_1(fifo_w_PE_3_5_V_V_full_n_pass_1_out),
    .PE_wrapper190_U0_fifo_w_out_V_V_write_pass_1(PE_wrapper190_U0_fifo_w_out_V_V_write_pass_1_in),
    .PE_wrapper179_U0_fifo_cin_out_V_V_din_pass_1(PE_wrapper179_U0_fifo_cin_out_V_V_din_pass_1_in),
    .fifo_cin_PE_3_5_V_V_full_n_pass_1(fifo_cin_PE_3_5_V_V_full_n_pass_1_out),
    .PE_wrapper179_U0_fifo_cin_out_V_V_write_pass_1(PE_wrapper179_U0_fifo_cin_out_V_V_write_pass_1_in),
    .PE_wrapper180_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper180_U0_fifo_cin_out_V_V_din_pass_0_in),
    .fifo_cin_PE_3_6_V_V_full_n_pass_0(fifo_cin_PE_3_6_V_V_full_n_pass_0_out),
    .PE_wrapper180_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper180_U0_fifo_cin_out_V_V_write_pass_0_in),
    .ap_clk(ap_clk),
    .ap_start_Boundary_X4Y6_To_X6Y6(ap_start_Boundary_X4Y6_To_X6Y6_in),
    .ap_rst_n_Boundary_X4Y6_To_X6Y6(ap_rst_n_Boundary_X4Y6_To_X6Y6_in),
    .ap_done_Boundary_X4Y6_To_X6Y6(ap_done_Boundary_X4Y6_To_X6Y6_out),
    .ap_start_Boundary_X4Y8_To_X6Y8(ap_start_Boundary_X4Y8_To_X6Y8_out),
    .ap_rst_n_Boundary_X4Y8_To_X6Y8(ap_rst_n_Boundary_X4Y8_To_X6Y8_out),
    .ap_done_Boundary_X4Y8_To_X6Y8(ap_done_Boundary_X4Y8_To_X6Y8_in)
  );


  (* keep_hierarchy = "yes" *) CR_X6Y4_To_CR_X7Y5_ctrl CR_X6Y4_To_CR_X7Y5_ctrl_U0 (
    .cout_drain_IO_L2_out568_U0_fifo_cout_drain_out_V_V_din_pass_1(cout_drain_IO_L2_out568_U0_fifo_cout_drain_out_V_V_din_pass_1_in),
    .cout_drain_IO_L2_out568_U0_fifo_cout_drain_out_V_V_din_pass_2(cout_drain_IO_L2_out568_U0_fifo_cout_drain_out_V_V_din_pass_2_out),
    .fifo_cout_drain_cout_drain_IO_L2_out_0_V_V_full_n_pass_1(fifo_cout_drain_cout_drain_IO_L2_out_0_V_V_full_n_pass_1_out),
    .fifo_cout_drain_cout_drain_IO_L2_out_0_V_V_full_n_pass_2(fifo_cout_drain_cout_drain_IO_L2_out_0_V_V_full_n_pass_2_in),
    .cout_drain_IO_L2_out568_U0_fifo_cout_drain_out_V_V_write_pass_1(cout_drain_IO_L2_out568_U0_fifo_cout_drain_out_V_V_write_pass_1_in),
    .cout_drain_IO_L2_out568_U0_fifo_cout_drain_out_V_V_write_pass_2(cout_drain_IO_L2_out568_U0_fifo_cout_drain_out_V_V_write_pass_2_out),
    .PE_wrapper165_U0_fifo_w_out_V_V_din_pass_1(PE_wrapper165_U0_fifo_w_out_V_V_din_pass_1_in),
    .fifo_w_PE_1_4_V_V_full_n_pass_1(fifo_w_PE_1_4_V_V_full_n_pass_1_out),
    .PE_wrapper165_U0_fifo_w_out_V_V_write_pass_1(PE_wrapper165_U0_fifo_w_out_V_V_write_pass_1_in),
    .cout_drain_IO_L2_out564_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L2_out564_U0_fifo_cout_drain_out_V_V_din_pass_0_out),
    .fifo_cout_drain_cout_drain_IO_L2_out_4_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L2_out_4_V_V_full_n_pass_0_in),
    .cout_drain_IO_L2_out564_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L2_out564_U0_fifo_cout_drain_out_V_V_write_pass_0_out),
    .cin_IO_L2_in127_U0_fifo_cin_out_V_V_din_pass_1(cin_IO_L2_in127_U0_fifo_cin_out_V_V_din_pass_1_in),
    .fifo_cin_cin_IO_L2_in_4_V_V_full_n_pass_1(fifo_cin_cin_IO_L2_in_4_V_V_full_n_pass_1_out),
    .cin_IO_L2_in127_U0_fifo_cin_out_V_V_write_pass_1(cin_IO_L2_in127_U0_fifo_cin_out_V_V_write_pass_1_in),
    .PE_wrapper179_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper179_U0_fifo_w_out_V_V_din_pass_0_out),
    .fifo_w_PE_2_6_V_V_full_n_pass_0(fifo_w_PE_2_6_V_V_full_n_pass_0_in),
    .PE_wrapper179_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper179_U0_fifo_w_out_V_V_write_pass_0_out),
    .cin_IO_L2_in128_U0_fifo_cin_out_V_V_din_pass_0(cin_IO_L2_in128_U0_fifo_cin_out_V_V_din_pass_0_out),
    .fifo_cin_cin_IO_L2_in_5_V_V_full_n_pass_0(fifo_cin_cin_IO_L2_in_5_V_V_full_n_pass_0_in),
    .cin_IO_L2_in128_U0_fifo_cin_out_V_V_write_pass_0(cin_IO_L2_in128_U0_fifo_cin_out_V_V_write_pass_0_out),
    .PE_wrapper179_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper179_U0_fifo_cout_drain_out_V_din_pass_0_out),
    .fifo_cout_drain_PE_2_5_V_full_n_pass_0(fifo_cout_drain_PE_2_5_V_full_n_pass_0_in),
    .PE_wrapper179_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper179_U0_fifo_cout_drain_out_V_write_pass_0_out),
    .PE_wrapper177_U0_fifo_w_out_V_V_din_pass_1(PE_wrapper177_U0_fifo_w_out_V_V_din_pass_1_in),
    .fifo_w_PE_2_4_V_V_full_n_pass_1(fifo_w_PE_2_4_V_V_full_n_pass_1_out),
    .PE_wrapper177_U0_fifo_w_out_V_V_write_pass_1(PE_wrapper177_U0_fifo_w_out_V_V_write_pass_1_in),
    .PE_wrapper153_U0_fifo_w_out_V_V_din_pass_1(PE_wrapper153_U0_fifo_w_out_V_V_din_pass_1_in),
    .fifo_w_PE_0_4_V_V_full_n_pass_1(fifo_w_PE_0_4_V_V_full_n_pass_1_out),
    .PE_wrapper153_U0_fifo_w_out_V_V_write_pass_1(PE_wrapper153_U0_fifo_w_out_V_V_write_pass_1_in),
    .PE_wrapper190_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper190_U0_fifo_cin_out_V_V_din_pass_0_out),
    .fifo_cin_PE_4_4_V_V_full_n_pass_0(fifo_cin_PE_4_4_V_V_full_n_pass_0_in),
    .PE_wrapper190_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper190_U0_fifo_cin_out_V_V_write_pass_0_out),
    .PE_wrapper166_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper166_U0_fifo_w_out_V_V_din_pass_0_out),
    .fifo_w_PE_1_5_V_V_full_n_pass_0(fifo_w_PE_1_5_V_V_full_n_pass_0_in),
    .PE_wrapper166_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper166_U0_fifo_w_out_V_V_write_pass_0_out),
    .PE_wrapper154_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper154_U0_fifo_w_out_V_V_din_pass_0_out),
    .fifo_w_PE_0_5_V_V_full_n_pass_0(fifo_w_PE_0_5_V_V_full_n_pass_0_in),
    .PE_wrapper154_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper154_U0_fifo_w_out_V_V_write_pass_0_out),
    .cout_drain_IO_L2_out563_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L2_out563_U0_fifo_cout_drain_out_V_V_din_pass_0_in),
    .fifo_cout_drain_cout_drain_IO_L2_out_5_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L2_out_5_V_V_full_n_pass_0_out),
    .cout_drain_IO_L2_out563_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L2_out563_U0_fifo_cout_drain_out_V_V_write_pass_0_in),
    .PE_wrapper190_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper190_U0_fifo_w_out_V_V_din_pass_0_out),
    .fifo_w_PE_3_5_V_V_full_n_pass_0(fifo_w_PE_3_5_V_V_full_n_pass_0_in),
    .PE_wrapper190_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper190_U0_fifo_w_out_V_V_write_pass_0_out),
    .PE_wrapper179_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper179_U0_fifo_cin_out_V_V_din_pass_0_out),
    .fifo_cin_PE_3_5_V_V_full_n_pass_0(fifo_cin_PE_3_5_V_V_full_n_pass_0_in),
    .PE_wrapper179_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper179_U0_fifo_cin_out_V_V_write_pass_0_out),
    .PE_wrapper202_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper202_U0_fifo_cout_drain_out_V_din_pass_0_in),
    .fifo_cout_drain_PE_4_4_V_full_n_pass_0(fifo_cout_drain_PE_4_4_V_full_n_pass_0_out),
    .PE_wrapper202_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper202_U0_fifo_cout_drain_out_V_write_pass_0_in),
    .PE_wrapper189_U0_fifo_w_out_V_V_din_pass_1(PE_wrapper189_U0_fifo_w_out_V_V_din_pass_1_in),
    .fifo_w_PE_3_4_V_V_full_n_pass_1(fifo_w_PE_3_4_V_V_full_n_pass_1_out),
    .PE_wrapper189_U0_fifo_w_out_V_V_write_pass_1(PE_wrapper189_U0_fifo_w_out_V_V_write_pass_1_in),
    .PE_wrapper167_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper167_U0_fifo_cin_out_V_V_din_pass_0_in),
    .fifo_cin_PE_2_5_V_V_full_n_pass_0(fifo_cin_PE_2_5_V_V_full_n_pass_0_out),
    .PE_wrapper167_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper167_U0_fifo_cin_out_V_V_write_pass_0_in),
    .cout_drain_IO_L1_out_wrapper441_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper441_U0_fifo_cout_drain_out_V_V_din_pass_0_in),
    .fifo_cout_drain_cout_drain_IO_L1_out_4_5_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_4_5_V_V_full_n_pass_0_out),
    .cout_drain_IO_L1_out_wrapper441_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper441_U0_fifo_cout_drain_out_V_V_write_pass_0_in),
    .ap_clk(ap_clk),
    .ap_start_Boundary_X6Y4_To_X8Y4(ap_start_Boundary_X6Y4_To_X8Y4_in),
    .ap_rst_n_Boundary_X6Y4_To_X8Y4(ap_rst_n_Boundary_X6Y4_To_X8Y4_in),
    .ap_done_Boundary_X6Y4_To_X8Y4(ap_done_Boundary_X6Y4_To_X8Y4_out),
    .ap_start_Boundary_X6Y6_To_X8Y6(ap_start_Boundary_X6Y6_To_X8Y6_out),
    .ap_rst_n_Boundary_X6Y6_To_X8Y6(ap_rst_n_Boundary_X6Y6_To_X8Y6_out),
    .ap_done_Boundary_X6Y6_To_X8Y6(ap_done_Boundary_X6Y6_To_X8Y6_in)
  );


  (* keep_hierarchy = "yes" *) CR_X6Y6_To_CR_X7Y7_ctrl CR_X6Y6_To_CR_X7Y7_ctrl_U0 (
    .PE_wrapper192_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper192_U0_fifo_w_out_V_V_din_pass_0_in),
    .PE_wrapper192_U0_fifo_w_out_V_V_din_pass_1(PE_wrapper192_U0_fifo_w_out_V_V_din_pass_1_out),
    .fifo_w_PE_3_7_V_V_full_n_pass_0(fifo_w_PE_3_7_V_V_full_n_pass_0_out),
    .fifo_w_PE_3_7_V_V_full_n_pass_1(fifo_w_PE_3_7_V_V_full_n_pass_1_in),
    .PE_wrapper192_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper192_U0_fifo_w_out_V_V_write_pass_0_in),
    .PE_wrapper192_U0_fifo_w_out_V_V_write_pass_1(PE_wrapper192_U0_fifo_w_out_V_V_write_pass_1_out),
    .cout_drain_IO_L2_out568_U0_fifo_cout_drain_out_V_V_din_pass_2(cout_drain_IO_L2_out568_U0_fifo_cout_drain_out_V_V_din_pass_2_in),
    .cout_drain_IO_L2_out568_U0_fifo_cout_drain_out_V_V_din_pass_3(cout_drain_IO_L2_out568_U0_fifo_cout_drain_out_V_V_din_pass_3_out),
    .fifo_cout_drain_cout_drain_IO_L2_out_0_V_V_full_n_pass_2(fifo_cout_drain_cout_drain_IO_L2_out_0_V_V_full_n_pass_2_out),
    .fifo_cout_drain_cout_drain_IO_L2_out_0_V_V_full_n_pass_3(fifo_cout_drain_cout_drain_IO_L2_out_0_V_V_full_n_pass_3_in),
    .cout_drain_IO_L2_out568_U0_fifo_cout_drain_out_V_V_write_pass_2(cout_drain_IO_L2_out568_U0_fifo_cout_drain_out_V_V_write_pass_2_in),
    .cout_drain_IO_L2_out568_U0_fifo_cout_drain_out_V_V_write_pass_3(cout_drain_IO_L2_out568_U0_fifo_cout_drain_out_V_V_write_pass_3_out),
    .PE_wrapper168_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper168_U0_fifo_w_out_V_V_din_pass_0_out),
    .fifo_w_PE_1_7_V_V_full_n_pass_0(fifo_w_PE_1_7_V_V_full_n_pass_0_in),
    .PE_wrapper168_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper168_U0_fifo_w_out_V_V_write_pass_0_out),
    .PE_wrapper179_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper179_U0_fifo_w_out_V_V_din_pass_0_in),
    .fifo_w_PE_2_6_V_V_full_n_pass_0(fifo_w_PE_2_6_V_V_full_n_pass_0_out),
    .PE_wrapper179_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper179_U0_fifo_w_out_V_V_write_pass_0_in),
    .cin_IO_L2_in128_U0_fifo_cin_out_V_V_din_pass_0(cin_IO_L2_in128_U0_fifo_cin_out_V_V_din_pass_0_in),
    .fifo_cin_cin_IO_L2_in_5_V_V_full_n_pass_0(fifo_cin_cin_IO_L2_in_5_V_V_full_n_pass_0_out),
    .cin_IO_L2_in128_U0_fifo_cin_out_V_V_write_pass_0(cin_IO_L2_in128_U0_fifo_cin_out_V_V_write_pass_0_in),
    .cout_drain_IO_L2_out561_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L2_out561_U0_fifo_cout_drain_out_V_V_din_pass_0_in),
    .fifo_cout_drain_cout_drain_IO_L2_out_7_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L2_out_7_V_V_full_n_pass_0_out),
    .cout_drain_IO_L2_out561_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L2_out561_U0_fifo_cout_drain_out_V_V_write_pass_0_in),
    .PE_wrapper242_U0_fifo_w_out_V_V_din_pass_2(PE_wrapper242_U0_fifo_w_out_V_V_din_pass_2_in),
    .fifo_w_PE_7_9_V_V_full_n_pass_2(fifo_w_PE_7_9_V_V_full_n_pass_2_out),
    .PE_wrapper242_U0_fifo_w_out_V_V_write_pass_2(PE_wrapper242_U0_fifo_w_out_V_V_write_pass_2_in),
    .PE_wrapper179_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper179_U0_fifo_cout_drain_out_V_din_pass_0_in),
    .fifo_cout_drain_PE_2_5_V_full_n_pass_0(fifo_cout_drain_PE_2_5_V_full_n_pass_0_out),
    .PE_wrapper179_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper179_U0_fifo_cout_drain_out_V_write_pass_0_in),
    .cin_IO_L2_in130_U0_fifo_cin_out_V_V_din_pass_0(cin_IO_L2_in130_U0_fifo_cin_out_V_V_din_pass_0_out),
    .fifo_cin_cin_IO_L2_in_7_V_V_full_n_pass_0(fifo_cin_cin_IO_L2_in_7_V_V_full_n_pass_0_in),
    .cin_IO_L2_in130_U0_fifo_cin_out_V_V_write_pass_0(cin_IO_L2_in130_U0_fifo_cin_out_V_V_write_pass_0_out),
    .PE_wrapper166_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper166_U0_fifo_w_out_V_V_din_pass_0_in),
    .fifo_w_PE_1_5_V_V_full_n_pass_0(fifo_w_PE_1_5_V_V_full_n_pass_0_out),
    .PE_wrapper166_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper166_U0_fifo_w_out_V_V_write_pass_0_in),
    .PE_wrapper243_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper243_U0_fifo_w_out_V_V_din_pass_0_out),
    .fifo_w_PE_7_10_V_V_full_n_pass_0(fifo_w_PE_7_10_V_V_full_n_pass_0_in),
    .PE_wrapper243_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper243_U0_fifo_w_out_V_V_write_pass_0_out),
    .PE_wrapper243_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper243_U0_fifo_cout_drain_out_V_din_pass_0_out),
    .fifo_cout_drain_PE_7_9_V_full_n_pass_0(fifo_cout_drain_PE_7_9_V_full_n_pass_0_in),
    .PE_wrapper243_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper243_U0_fifo_cout_drain_out_V_write_pass_0_out),
    .PE_wrapper243_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper243_U0_fifo_cin_out_V_V_din_pass_0_out),
    .fifo_cin_PE_8_9_V_V_full_n_pass_0(fifo_cin_PE_8_9_V_V_full_n_pass_0_in),
    .PE_wrapper243_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper243_U0_fifo_cin_out_V_V_write_pass_0_out),
    .PE_wrapper154_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper154_U0_fifo_w_out_V_V_din_pass_0_in),
    .fifo_w_PE_0_5_V_V_full_n_pass_0(fifo_w_PE_0_5_V_V_full_n_pass_0_out),
    .PE_wrapper154_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper154_U0_fifo_w_out_V_V_write_pass_0_in),
    .PE_wrapper156_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper156_U0_fifo_w_out_V_V_din_pass_0_out),
    .fifo_w_PE_0_7_V_V_full_n_pass_0(fifo_w_PE_0_7_V_V_full_n_pass_0_in),
    .PE_wrapper156_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper156_U0_fifo_w_out_V_V_write_pass_0_out),
    .PE_wrapper180_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper180_U0_fifo_cin_out_V_V_din_pass_0_out),
    .fifo_cin_PE_3_6_V_V_full_n_pass_0(fifo_cin_PE_3_6_V_V_full_n_pass_0_in),
    .PE_wrapper180_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper180_U0_fifo_cin_out_V_V_write_pass_0_out),
    .cout_drain_IO_L2_out563_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L2_out563_U0_fifo_cout_drain_out_V_V_din_pass_0_out),
    .fifo_cout_drain_cout_drain_IO_L2_out_5_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L2_out_5_V_V_full_n_pass_0_in),
    .cout_drain_IO_L2_out563_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L2_out563_U0_fifo_cout_drain_out_V_V_write_pass_0_out),
    .PE_wrapper191_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper191_U0_fifo_cout_drain_out_V_din_pass_0_in),
    .fifo_cout_drain_PE_3_5_V_full_n_pass_0(fifo_cout_drain_PE_3_5_V_full_n_pass_0_out),
    .PE_wrapper191_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper191_U0_fifo_cout_drain_out_V_write_pass_0_in),
    .cout_drain_IO_L1_out_wrapper474_U0_fifo_cout_drain_out_V_V_din_pass_1(cout_drain_IO_L1_out_wrapper474_U0_fifo_cout_drain_out_V_V_din_pass_1_in),
    .fifo_cout_drain_cout_drain_IO_L1_out_6_4_V_V_full_n_pass_1(fifo_cout_drain_cout_drain_IO_L1_out_6_4_V_V_full_n_pass_1_out),
    .cout_drain_IO_L1_out_wrapper474_U0_fifo_cout_drain_out_V_V_write_pass_1(cout_drain_IO_L1_out_wrapper474_U0_fifo_cout_drain_out_V_V_write_pass_1_in),
    .cout_drain_IO_L1_out_wrapper458_U0_fifo_cout_drain_out_V_V_din_pass_1(cout_drain_IO_L1_out_wrapper458_U0_fifo_cout_drain_out_V_V_din_pass_1_in),
    .fifo_cout_drain_cout_drain_IO_L1_out_5_4_V_V_full_n_pass_1(fifo_cout_drain_cout_drain_IO_L1_out_5_4_V_V_full_n_pass_1_out),
    .cout_drain_IO_L1_out_wrapper458_U0_fifo_cout_drain_out_V_V_write_pass_1(cout_drain_IO_L1_out_wrapper458_U0_fifo_cout_drain_out_V_V_write_pass_1_in),
    .PE_wrapper180_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper180_U0_fifo_w_out_V_V_din_pass_0_out),
    .fifo_w_PE_2_7_V_V_full_n_pass_0(fifo_w_PE_2_7_V_V_full_n_pass_0_in),
    .PE_wrapper180_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper180_U0_fifo_w_out_V_V_write_pass_0_out),
    .PE_wrapper167_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper167_U0_fifo_cin_out_V_V_din_pass_0_out),
    .fifo_cin_PE_2_5_V_V_full_n_pass_0(fifo_cin_PE_2_5_V_V_full_n_pass_0_in),
    .PE_wrapper167_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper167_U0_fifo_cin_out_V_V_write_pass_0_out),
    .PE_wrapper192_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper192_U0_fifo_cout_drain_out_V_din_pass_0_in),
    .fifo_cout_drain_PE_3_6_V_full_n_pass_0(fifo_cout_drain_PE_3_6_V_full_n_pass_0_out),
    .PE_wrapper192_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper192_U0_fifo_cout_drain_out_V_write_pass_0_in),
    .PE_wrapper231_U0_fifo_cin_out_V_V_din_pass_4(PE_wrapper231_U0_fifo_cin_out_V_V_din_pass_4_in),
    .fifo_cin_PE_7_9_V_V_full_n_pass_4(fifo_cin_PE_7_9_V_V_full_n_pass_4_out),
    .PE_wrapper231_U0_fifo_cin_out_V_V_write_pass_4(PE_wrapper231_U0_fifo_cin_out_V_V_write_pass_4_in),
    .ap_clk(ap_clk),
    .ap_start_Boundary_X6Y6_To_X8Y6(ap_start_Boundary_X6Y6_To_X8Y6_in),
    .ap_rst_n_Boundary_X6Y6_To_X8Y6(ap_rst_n_Boundary_X6Y6_To_X8Y6_in),
    .ap_done_Boundary_X6Y6_To_X8Y6(ap_done_Boundary_X6Y6_To_X8Y6_out),
    .ap_start_Boundary_X6Y8_To_X8Y8(ap_start_Boundary_X6Y8_To_X8Y8_out),
    .ap_rst_n_Boundary_X6Y8_To_X8Y8(ap_rst_n_Boundary_X6Y8_To_X8Y8_out),
    .ap_done_Boundary_X6Y8_To_X8Y8(ap_done_Boundary_X6Y8_To_X8Y8_in)
  );


  (* keep_hierarchy = "yes" *) CR_X4Y8_To_CR_X5Y9_ctrl CR_X4Y8_To_CR_X5Y9_ctrl_U0 (
    .PE_wrapper251_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper251_U0_fifo_w_out_V_V_din_pass_0_in),
    .PE_wrapper251_U0_fifo_w_out_V_V_din_pass_1(PE_wrapper251_U0_fifo_w_out_V_V_din_pass_1_out),
    .fifo_w_PE_8_6_V_V_full_n_pass_0(fifo_w_PE_8_6_V_V_full_n_pass_0_out),
    .fifo_w_PE_8_6_V_V_full_n_pass_1(fifo_w_PE_8_6_V_V_full_n_pass_1_in),
    .PE_wrapper251_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper251_U0_fifo_w_out_V_V_write_pass_0_in),
    .PE_wrapper251_U0_fifo_w_out_V_V_write_pass_1(PE_wrapper251_U0_fifo_w_out_V_V_write_pass_1_out),
    .PE_wrapper239_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper239_U0_fifo_w_out_V_V_din_pass_0_in),
    .PE_wrapper239_U0_fifo_w_out_V_V_din_pass_1(PE_wrapper239_U0_fifo_w_out_V_V_din_pass_1_out),
    .fifo_w_PE_7_6_V_V_full_n_pass_0(fifo_w_PE_7_6_V_V_full_n_pass_0_out),
    .fifo_w_PE_7_6_V_V_full_n_pass_1(fifo_w_PE_7_6_V_V_full_n_pass_1_in),
    .PE_wrapper239_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper239_U0_fifo_w_out_V_V_write_pass_0_in),
    .PE_wrapper239_U0_fifo_w_out_V_V_write_pass_1(PE_wrapper239_U0_fifo_w_out_V_V_write_pass_1_out),
    .cout_drain_IO_L1_out_wrapper469_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper469_U0_fifo_cout_drain_out_V_V_din_pass_0_in),
    .cout_drain_IO_L1_out_wrapper469_U0_fifo_cout_drain_out_V_V_din_pass_1(cout_drain_IO_L1_out_wrapper469_U0_fifo_cout_drain_out_V_V_din_pass_1_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_6_9_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_6_9_V_V_full_n_pass_0_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_6_9_V_V_full_n_pass_1(fifo_cout_drain_cout_drain_IO_L1_out_6_9_V_V_full_n_pass_1_in),
    .cout_drain_IO_L1_out_wrapper469_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper469_U0_fifo_cout_drain_out_V_V_write_pass_0_in),
    .cout_drain_IO_L1_out_wrapper469_U0_fifo_cout_drain_out_V_V_write_pass_1(cout_drain_IO_L1_out_wrapper469_U0_fifo_cout_drain_out_V_V_write_pass_1_out),
    .kernel0_entry12_U0_cout_V_out_din_pass_3(kernel0_entry12_U0_cout_V_out_din_pass_3_in),
    .kernel0_entry12_U0_cout_V_out_din_pass_4(kernel0_entry12_U0_cout_V_out_din_pass_4_out),
    .cout_V_c_full_n_pass_3(cout_V_c_full_n_pass_3_out),
    .cout_V_c_full_n_pass_4(cout_V_c_full_n_pass_4_in),
    .kernel0_entry12_U0_cout_V_out_write_pass_3(kernel0_entry12_U0_cout_V_out_write_pass_3_in),
    .kernel0_entry12_U0_cout_V_out_write_pass_4(kernel0_entry12_U0_cout_V_out_write_pass_4_out),
    .PE_wrapper243_U0_fifo_w_out_V_V_din_pass_1(PE_wrapper243_U0_fifo_w_out_V_V_din_pass_1_in),
    .PE_wrapper243_U0_fifo_w_out_V_V_din_pass_2(PE_wrapper243_U0_fifo_w_out_V_V_din_pass_2_out),
    .fifo_w_PE_7_10_V_V_full_n_pass_1(fifo_w_PE_7_10_V_V_full_n_pass_1_out),
    .fifo_w_PE_7_10_V_V_full_n_pass_2(fifo_w_PE_7_10_V_V_full_n_pass_2_in),
    .PE_wrapper243_U0_fifo_w_out_V_V_write_pass_1(PE_wrapper243_U0_fifo_w_out_V_V_write_pass_1_in),
    .PE_wrapper243_U0_fifo_w_out_V_V_write_pass_2(PE_wrapper243_U0_fifo_w_out_V_V_write_pass_2_out),
    .PE_wrapper243_U0_fifo_cout_drain_out_V_din_pass_1(PE_wrapper243_U0_fifo_cout_drain_out_V_din_pass_1_in),
    .PE_wrapper243_U0_fifo_cout_drain_out_V_din_pass_2(PE_wrapper243_U0_fifo_cout_drain_out_V_din_pass_2_out),
    .fifo_cout_drain_PE_7_9_V_full_n_pass_1(fifo_cout_drain_PE_7_9_V_full_n_pass_1_out),
    .fifo_cout_drain_PE_7_9_V_full_n_pass_2(fifo_cout_drain_PE_7_9_V_full_n_pass_2_in),
    .PE_wrapper243_U0_fifo_cout_drain_out_V_write_pass_1(PE_wrapper243_U0_fifo_cout_drain_out_V_write_pass_1_in),
    .PE_wrapper243_U0_fifo_cout_drain_out_V_write_pass_2(PE_wrapper243_U0_fifo_cout_drain_out_V_write_pass_2_out),
    .PE_wrapper243_U0_fifo_cin_out_V_V_din_pass_1(PE_wrapper243_U0_fifo_cin_out_V_V_din_pass_1_in),
    .PE_wrapper243_U0_fifo_cin_out_V_V_din_pass_2(PE_wrapper243_U0_fifo_cin_out_V_V_din_pass_2_out),
    .fifo_cin_PE_8_9_V_V_full_n_pass_1(fifo_cin_PE_8_9_V_V_full_n_pass_1_out),
    .fifo_cin_PE_8_9_V_V_full_n_pass_2(fifo_cin_PE_8_9_V_V_full_n_pass_2_in),
    .PE_wrapper243_U0_fifo_cin_out_V_V_write_pass_1(PE_wrapper243_U0_fifo_cin_out_V_V_write_pass_1_in),
    .PE_wrapper243_U0_fifo_cin_out_V_V_write_pass_2(PE_wrapper243_U0_fifo_cin_out_V_V_write_pass_2_out),
    .cout_drain_IO_L3_out_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L3_out_U0_fifo_cout_drain_out_V_V_din_pass_0_in),
    .cout_drain_IO_L3_out_U0_fifo_cout_drain_out_V_V_din_pass_1(cout_drain_IO_L3_out_U0_fifo_cout_drain_out_V_V_din_pass_1_out),
    .fifo_cout_drain_cout_drain_IO_L3_out_serialize_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L3_out_serialize_V_V_full_n_pass_0_out),
    .fifo_cout_drain_cout_drain_IO_L3_out_serialize_V_V_full_n_pass_1(fifo_cout_drain_cout_drain_IO_L3_out_serialize_V_V_full_n_pass_1_in),
    .cout_drain_IO_L3_out_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L3_out_U0_fifo_cout_drain_out_V_V_write_pass_0_in),
    .cout_drain_IO_L3_out_U0_fifo_cout_drain_out_V_V_write_pass_1(cout_drain_IO_L3_out_U0_fifo_cout_drain_out_V_V_write_pass_1_out),
    .PE_wrapper192_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper192_U0_fifo_cin_out_V_V_din_pass_0_in),
    .fifo_cin_PE_4_6_V_V_full_n_pass_0(fifo_cin_PE_4_6_V_V_full_n_pass_0_out),
    .PE_wrapper192_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper192_U0_fifo_cin_out_V_V_write_pass_0_in),
    .cout_drain_IO_L1_out_wrapper471_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper471_U0_fifo_cout_drain_out_V_V_din_pass_0_in),
    .fifo_cout_drain_cout_drain_IO_L1_out_6_7_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_6_7_V_V_full_n_pass_0_out),
    .cout_drain_IO_L1_out_wrapper471_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper471_U0_fifo_cout_drain_out_V_V_write_pass_0_in),
    .PE_wrapper214_U0_fifo_w_out_V_V_din_pass_1(PE_wrapper214_U0_fifo_w_out_V_V_din_pass_1_in),
    .fifo_w_PE_5_5_V_V_full_n_pass_1(fifo_w_PE_5_5_V_V_full_n_pass_1_out),
    .PE_wrapper214_U0_fifo_w_out_V_V_write_pass_1(PE_wrapper214_U0_fifo_w_out_V_V_write_pass_1_in),
    .cout_drain_IO_L1_out_wrapper490_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper490_U0_fifo_cout_drain_out_V_V_din_pass_0_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_7_4_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_7_4_V_V_full_n_pass_0_in),
    .cout_drain_IO_L1_out_wrapper490_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper490_U0_fifo_cout_drain_out_V_V_write_pass_0_out),
    .PE_wrapper205_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper205_U0_fifo_cin_out_V_V_din_pass_0_in),
    .fifo_cin_PE_5_7_V_V_full_n_pass_0(fifo_cin_PE_5_7_V_V_full_n_pass_0_out),
    .PE_wrapper205_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper205_U0_fifo_cin_out_V_V_write_pass_0_in),
    .PE_wrapper217_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper217_U0_fifo_w_out_V_V_din_pass_0_out),
    .fifo_w_PE_5_8_V_V_full_n_pass_0(fifo_w_PE_5_8_V_V_full_n_pass_0_in),
    .PE_wrapper217_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper217_U0_fifo_w_out_V_V_write_pass_0_out),
    .PE_wrapper215_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper215_U0_fifo_cin_out_V_V_din_pass_0_out),
    .fifo_cin_PE_6_5_V_V_full_n_pass_0(fifo_cin_PE_6_5_V_V_full_n_pass_0_in),
    .PE_wrapper215_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper215_U0_fifo_cin_out_V_V_write_pass_0_out),
    .PE_wrapper227_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper227_U0_fifo_w_out_V_V_din_pass_0_in),
    .fifo_w_PE_6_6_V_V_full_n_pass_0(fifo_w_PE_6_6_V_V_full_n_pass_0_out),
    .PE_wrapper227_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper227_U0_fifo_w_out_V_V_write_pass_0_in),
    .PE_wrapper228_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper228_U0_fifo_cin_out_V_V_din_pass_0_out),
    .fifo_cin_PE_7_6_V_V_full_n_pass_0(fifo_cin_PE_7_6_V_V_full_n_pass_0_in),
    .PE_wrapper228_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper228_U0_fifo_cin_out_V_V_write_pass_0_out),
    .cout_drain_IO_L1_out_wrapper474_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper474_U0_fifo_cout_drain_out_V_V_din_pass_0_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_6_4_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_6_4_V_V_full_n_pass_0_in),
    .cout_drain_IO_L1_out_wrapper474_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper474_U0_fifo_cout_drain_out_V_V_write_pass_0_out),
    .cout_drain_IO_L1_out_wrapper458_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper458_U0_fifo_cout_drain_out_V_V_din_pass_0_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_5_4_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_5_4_V_V_full_n_pass_0_in),
    .cout_drain_IO_L1_out_wrapper458_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper458_U0_fifo_cout_drain_out_V_V_write_pass_0_out),
    .PE_wrapper229_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper229_U0_fifo_w_out_V_V_din_pass_0_out),
    .fifo_w_PE_6_8_V_V_full_n_pass_0(fifo_w_PE_6_8_V_V_full_n_pass_0_in),
    .PE_wrapper229_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper229_U0_fifo_w_out_V_V_write_pass_0_out),
    .PE_wrapper202_U0_fifo_w_out_V_V_din_pass_1(PE_wrapper202_U0_fifo_w_out_V_V_din_pass_1_in),
    .fifo_w_PE_4_5_V_V_full_n_pass_1(fifo_w_PE_4_5_V_V_full_n_pass_1_out),
    .PE_wrapper202_U0_fifo_w_out_V_V_write_pass_1(PE_wrapper202_U0_fifo_w_out_V_V_write_pass_1_in),
    .cout_drain_IO_L1_out_wrapper456_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper456_U0_fifo_cout_drain_out_V_V_din_pass_0_in),
    .fifo_cout_drain_cout_drain_IO_L1_out_5_6_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_5_6_V_V_full_n_pass_0_out),
    .cout_drain_IO_L1_out_wrapper456_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper456_U0_fifo_cout_drain_out_V_V_write_pass_0_in),
    .PE_wrapper229_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper229_U0_fifo_cin_out_V_V_din_pass_0_out),
    .fifo_cin_PE_7_7_V_V_full_n_pass_0(fifo_cin_PE_7_7_V_V_full_n_pass_0_in),
    .PE_wrapper229_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper229_U0_fifo_cin_out_V_V_write_pass_0_out),
    .PE_wrapper191_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper191_U0_fifo_cin_out_V_V_din_pass_0_in),
    .fifo_cin_PE_4_5_V_V_full_n_pass_0(fifo_cin_PE_4_5_V_V_full_n_pass_0_out),
    .PE_wrapper191_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper191_U0_fifo_cin_out_V_V_write_pass_0_in),
    .PE_wrapper205_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper205_U0_fifo_cout_drain_out_V_din_pass_0_in),
    .fifo_cout_drain_PE_4_7_V_full_n_pass_0(fifo_cout_drain_PE_4_7_V_full_n_pass_0_out),
    .PE_wrapper205_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper205_U0_fifo_cout_drain_out_V_write_pass_0_in),
    .PE_wrapper204_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper204_U0_fifo_w_out_V_V_din_pass_0_out),
    .fifo_w_PE_4_7_V_V_full_n_pass_0(fifo_w_PE_4_7_V_V_full_n_pass_0_in),
    .PE_wrapper204_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper204_U0_fifo_w_out_V_V_write_pass_0_out),
    .cout_drain_IO_L1_out_wrapper487_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper487_U0_fifo_cout_drain_out_V_V_din_pass_0_in),
    .fifo_cout_drain_cout_drain_IO_L1_out_7_7_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_7_7_V_V_full_n_pass_0_out),
    .cout_drain_IO_L1_out_wrapper487_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper487_U0_fifo_cout_drain_out_V_V_write_pass_0_in),
    .ap_clk(ap_clk),
    .ap_start_Boundary_X4Y8_To_X6Y8(ap_start_Boundary_X4Y8_To_X6Y8_in),
    .ap_rst_n_Boundary_X4Y8_To_X6Y8(ap_rst_n_Boundary_X4Y8_To_X6Y8_in),
    .ap_done_Boundary_X4Y8_To_X6Y8(ap_done_Boundary_X4Y8_To_X6Y8_out),
    .ap_start_Boundary_X4Y10_To_X6Y10(ap_start_Boundary_X4Y10_To_X6Y10_out),
    .ap_rst_n_Boundary_X4Y10_To_X6Y10(ap_rst_n_Boundary_X4Y10_To_X6Y10_out),
    .ap_done_Boundary_X4Y10_To_X6Y10(ap_done_Boundary_X4Y10_To_X6Y10_in)
  );


  (* keep_hierarchy = "yes" *) CR_X4Y10_To_CR_X5Y11_ctrl CR_X4Y10_To_CR_X5Y11_ctrl_U0 (
    .kernel0_entry12_U0_cout_V_out_din_pass_4(kernel0_entry12_U0_cout_V_out_din_pass_4_in),
    .kernel0_entry12_U0_cout_V_out_din_pass_5(kernel0_entry12_U0_cout_V_out_din_pass_5_out),
    .cout_V_c_full_n_pass_4(cout_V_c_full_n_pass_4_out),
    .cout_V_c_full_n_pass_5(cout_V_c_full_n_pass_5_in),
    .kernel0_entry12_U0_cout_V_out_write_pass_4(kernel0_entry12_U0_cout_V_out_write_pass_4_in),
    .kernel0_entry12_U0_cout_V_out_write_pass_5(kernel0_entry12_U0_cout_V_out_write_pass_5_out),
    .PE_wrapper243_U0_fifo_w_out_V_V_din_pass_2(PE_wrapper243_U0_fifo_w_out_V_V_din_pass_2_in),
    .PE_wrapper243_U0_fifo_w_out_V_V_din_pass_3(PE_wrapper243_U0_fifo_w_out_V_V_din_pass_3_out),
    .fifo_w_PE_7_10_V_V_full_n_pass_2(fifo_w_PE_7_10_V_V_full_n_pass_2_out),
    .fifo_w_PE_7_10_V_V_full_n_pass_3(fifo_w_PE_7_10_V_V_full_n_pass_3_in),
    .PE_wrapper243_U0_fifo_w_out_V_V_write_pass_2(PE_wrapper243_U0_fifo_w_out_V_V_write_pass_2_in),
    .PE_wrapper243_U0_fifo_w_out_V_V_write_pass_3(PE_wrapper243_U0_fifo_w_out_V_V_write_pass_3_out),
    .PE_wrapper243_U0_fifo_cout_drain_out_V_din_pass_2(PE_wrapper243_U0_fifo_cout_drain_out_V_din_pass_2_in),
    .PE_wrapper243_U0_fifo_cout_drain_out_V_din_pass_3(PE_wrapper243_U0_fifo_cout_drain_out_V_din_pass_3_out),
    .fifo_cout_drain_PE_7_9_V_full_n_pass_2(fifo_cout_drain_PE_7_9_V_full_n_pass_2_out),
    .fifo_cout_drain_PE_7_9_V_full_n_pass_3(fifo_cout_drain_PE_7_9_V_full_n_pass_3_in),
    .PE_wrapper243_U0_fifo_cout_drain_out_V_write_pass_2(PE_wrapper243_U0_fifo_cout_drain_out_V_write_pass_2_in),
    .PE_wrapper243_U0_fifo_cout_drain_out_V_write_pass_3(PE_wrapper243_U0_fifo_cout_drain_out_V_write_pass_3_out),
    .PE_wrapper243_U0_fifo_cin_out_V_V_din_pass_2(PE_wrapper243_U0_fifo_cin_out_V_V_din_pass_2_in),
    .PE_wrapper243_U0_fifo_cin_out_V_V_din_pass_3(PE_wrapper243_U0_fifo_cin_out_V_V_din_pass_3_out),
    .fifo_cin_PE_8_9_V_V_full_n_pass_2(fifo_cin_PE_8_9_V_V_full_n_pass_2_out),
    .fifo_cin_PE_8_9_V_V_full_n_pass_3(fifo_cin_PE_8_9_V_V_full_n_pass_3_in),
    .PE_wrapper243_U0_fifo_cin_out_V_V_write_pass_2(PE_wrapper243_U0_fifo_cin_out_V_V_write_pass_2_in),
    .PE_wrapper243_U0_fifo_cin_out_V_V_write_pass_3(PE_wrapper243_U0_fifo_cin_out_V_V_write_pass_3_out),
    .PE_wrapper182_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper182_U0_fifo_w_out_V_V_din_pass_0_in),
    .PE_wrapper182_U0_fifo_w_out_V_V_din_pass_1(PE_wrapper182_U0_fifo_w_out_V_V_din_pass_1_out),
    .fifo_w_PE_2_9_V_V_full_n_pass_0(fifo_w_PE_2_9_V_V_full_n_pass_0_out),
    .fifo_w_PE_2_9_V_V_full_n_pass_1(fifo_w_PE_2_9_V_V_full_n_pass_1_in),
    .PE_wrapper182_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper182_U0_fifo_w_out_V_V_write_pass_0_in),
    .PE_wrapper182_U0_fifo_w_out_V_V_write_pass_1(PE_wrapper182_U0_fifo_w_out_V_V_write_pass_1_out),
    .cout_drain_IO_L3_out_U0_fifo_cout_drain_out_V_V_din_pass_1(cout_drain_IO_L3_out_U0_fifo_cout_drain_out_V_V_din_pass_1_in),
    .cout_drain_IO_L3_out_U0_fifo_cout_drain_out_V_V_din_pass_2(cout_drain_IO_L3_out_U0_fifo_cout_drain_out_V_V_din_pass_2_out),
    .fifo_cout_drain_cout_drain_IO_L3_out_serialize_V_V_full_n_pass_1(fifo_cout_drain_cout_drain_IO_L3_out_serialize_V_V_full_n_pass_1_out),
    .fifo_cout_drain_cout_drain_IO_L3_out_serialize_V_V_full_n_pass_2(fifo_cout_drain_cout_drain_IO_L3_out_serialize_V_V_full_n_pass_2_in),
    .cout_drain_IO_L3_out_U0_fifo_cout_drain_out_V_V_write_pass_1(cout_drain_IO_L3_out_U0_fifo_cout_drain_out_V_V_write_pass_1_in),
    .cout_drain_IO_L3_out_U0_fifo_cout_drain_out_V_V_write_pass_2(cout_drain_IO_L3_out_U0_fifo_cout_drain_out_V_V_write_pass_2_out),
    .PE_wrapper194_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper194_U0_fifo_w_out_V_V_din_pass_0_in),
    .PE_wrapper194_U0_fifo_w_out_V_V_din_pass_1(PE_wrapper194_U0_fifo_w_out_V_V_din_pass_1_out),
    .fifo_w_PE_3_9_V_V_full_n_pass_0(fifo_w_PE_3_9_V_V_full_n_pass_0_out),
    .fifo_w_PE_3_9_V_V_full_n_pass_1(fifo_w_PE_3_9_V_V_full_n_pass_1_in),
    .PE_wrapper194_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper194_U0_fifo_w_out_V_V_write_pass_0_in),
    .PE_wrapper194_U0_fifo_w_out_V_V_write_pass_1(PE_wrapper194_U0_fifo_w_out_V_V_write_pass_1_out),
    .PE_wrapper253_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper253_U0_fifo_cin_out_V_V_din_pass_0_out),
    .fifo_cin_PE_9_7_V_V_full_n_pass_0(fifo_cin_PE_9_7_V_V_full_n_pass_0_in),
    .PE_wrapper253_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper253_U0_fifo_cin_out_V_V_write_pass_0_out),
    .cout_drain_IO_L1_out_wrapper471_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper471_U0_fifo_cout_drain_out_V_V_din_pass_0_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_6_7_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_6_7_V_V_full_n_pass_0_in),
    .cout_drain_IO_L1_out_wrapper471_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper471_U0_fifo_cout_drain_out_V_V_write_pass_0_out),
    .PE_wrapper218_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper218_U0_fifo_cout_drain_out_V_din_pass_0_in),
    .fifo_cout_drain_PE_5_8_V_full_n_pass_0(fifo_cout_drain_PE_5_8_V_full_n_pass_0_out),
    .PE_wrapper218_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper218_U0_fifo_cout_drain_out_V_write_pass_0_in),
    .PE_wrapper242_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper242_U0_fifo_w_out_V_V_din_pass_0_out),
    .fifo_w_PE_7_9_V_V_full_n_pass_0(fifo_w_PE_7_9_V_V_full_n_pass_0_in),
    .PE_wrapper242_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper242_U0_fifo_w_out_V_V_write_pass_0_out),
    .PE_wrapper230_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper230_U0_fifo_w_out_V_V_din_pass_0_out),
    .fifo_w_PE_6_9_V_V_full_n_pass_0(fifo_w_PE_6_9_V_V_full_n_pass_0_in),
    .PE_wrapper230_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper230_U0_fifo_w_out_V_V_write_pass_0_out),
    .cout_drain_IO_L1_out_wrapper506_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper506_U0_fifo_cout_drain_out_V_V_din_pass_0_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_8_4_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_8_4_V_V_full_n_pass_0_in),
    .cout_drain_IO_L1_out_wrapper506_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper506_U0_fifo_cout_drain_out_V_V_write_pass_0_out),
    .PE_wrapper252_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper252_U0_fifo_cin_out_V_V_din_pass_0_out),
    .fifo_cin_PE_9_6_V_V_full_n_pass_0(fifo_cin_PE_9_6_V_V_full_n_pass_0_in),
    .PE_wrapper252_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper252_U0_fifo_cin_out_V_V_write_pass_0_out),
    .PE_wrapper228_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper228_U0_fifo_cin_out_V_V_din_pass_0_in),
    .fifo_cin_PE_7_6_V_V_full_n_pass_0(fifo_cin_PE_7_6_V_V_full_n_pass_0_out),
    .PE_wrapper228_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper228_U0_fifo_cin_out_V_V_write_pass_0_in),
    .PE_wrapper254_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper254_U0_fifo_w_out_V_V_din_pass_0_out),
    .fifo_w_PE_8_9_V_V_full_n_pass_0(fifo_w_PE_8_9_V_V_full_n_pass_0_in),
    .PE_wrapper254_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper254_U0_fifo_w_out_V_V_write_pass_0_out),
    .cout_drain_IO_L1_out_wrapper501_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper501_U0_fifo_cout_drain_out_V_V_din_pass_0_in),
    .fifo_cout_drain_cout_drain_IO_L1_out_8_9_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_8_9_V_V_full_n_pass_0_out),
    .cout_drain_IO_L1_out_wrapper501_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper501_U0_fifo_cout_drain_out_V_V_write_pass_0_in),
    .PE_wrapper229_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper229_U0_fifo_w_out_V_V_din_pass_0_in),
    .fifo_w_PE_6_8_V_V_full_n_pass_0(fifo_w_PE_6_8_V_V_full_n_pass_0_out),
    .PE_wrapper229_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper229_U0_fifo_w_out_V_V_write_pass_0_in),
    .PE_wrapper229_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper229_U0_fifo_cin_out_V_V_din_pass_0_in),
    .fifo_cin_PE_7_7_V_V_full_n_pass_0(fifo_cin_PE_7_7_V_V_full_n_pass_0_out),
    .PE_wrapper229_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper229_U0_fifo_cin_out_V_V_write_pass_0_in),
    .PE_wrapper251_U0_fifo_w_out_V_V_din_pass_1(PE_wrapper251_U0_fifo_w_out_V_V_din_pass_1_in),
    .fifo_w_PE_8_6_V_V_full_n_pass_1(fifo_w_PE_8_6_V_V_full_n_pass_1_out),
    .PE_wrapper251_U0_fifo_w_out_V_V_write_pass_1(PE_wrapper251_U0_fifo_w_out_V_V_write_pass_1_in),
    .cout_drain_IO_L1_out_wrapper485_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper485_U0_fifo_cout_drain_out_V_V_din_pass_0_in),
    .fifo_cout_drain_cout_drain_IO_L1_out_7_9_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_7_9_V_V_full_n_pass_0_out),
    .cout_drain_IO_L1_out_wrapper485_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper485_U0_fifo_cout_drain_out_V_V_write_pass_0_in),
    .cout_drain_IO_L1_out_wrapper487_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper487_U0_fifo_cout_drain_out_V_V_din_pass_0_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_7_7_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_7_7_V_V_full_n_pass_0_in),
    .cout_drain_IO_L1_out_wrapper487_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper487_U0_fifo_cout_drain_out_V_V_write_pass_0_out),
    .PE_wrapper206_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper206_U0_fifo_cout_drain_out_V_din_pass_0_in),
    .fifo_cout_drain_PE_4_8_V_full_n_pass_0(fifo_cout_drain_PE_4_8_V_full_n_pass_0_out),
    .PE_wrapper206_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper206_U0_fifo_cout_drain_out_V_write_pass_0_in),
    .PE_wrapper218_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper218_U0_fifo_cin_out_V_V_din_pass_0_in),
    .fifo_cin_PE_6_8_V_V_full_n_pass_0(fifo_cin_PE_6_8_V_V_full_n_pass_0_out),
    .PE_wrapper218_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper218_U0_fifo_cin_out_V_V_write_pass_0_in),
    .PE_wrapper239_U0_fifo_w_out_V_V_din_pass_1(PE_wrapper239_U0_fifo_w_out_V_V_din_pass_1_in),
    .fifo_w_PE_7_6_V_V_full_n_pass_1(fifo_w_PE_7_6_V_V_full_n_pass_1_out),
    .PE_wrapper239_U0_fifo_w_out_V_V_write_pass_1(PE_wrapper239_U0_fifo_w_out_V_V_write_pass_1_in),
    .PE_wrapper254_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper254_U0_fifo_cin_out_V_V_din_pass_0_out),
    .fifo_cin_PE_9_8_V_V_full_n_pass_0(fifo_cin_PE_9_8_V_V_full_n_pass_0_in),
    .PE_wrapper254_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper254_U0_fifo_cin_out_V_V_write_pass_0_out),
    .cout_drain_IO_L1_out_wrapper469_U0_fifo_cout_drain_out_V_V_din_pass_1(cout_drain_IO_L1_out_wrapper469_U0_fifo_cout_drain_out_V_V_din_pass_1_in),
    .fifo_cout_drain_cout_drain_IO_L1_out_6_9_V_V_full_n_pass_1(fifo_cout_drain_cout_drain_IO_L1_out_6_9_V_V_full_n_pass_1_out),
    .cout_drain_IO_L1_out_wrapper469_U0_fifo_cout_drain_out_V_V_write_pass_1(cout_drain_IO_L1_out_wrapper469_U0_fifo_cout_drain_out_V_V_write_pass_1_in),
    .ap_clk(ap_clk),
    .ap_start_Boundary_X4Y10_To_X6Y10(ap_start_Boundary_X4Y10_To_X6Y10_in),
    .ap_rst_n_Boundary_X4Y10_To_X6Y10(ap_rst_n_Boundary_X4Y10_To_X6Y10_in),
    .ap_done_Boundary_X4Y10_To_X6Y10(ap_done_Boundary_X4Y10_To_X6Y10_out),
    .ap_start_Boundary_X4Y12_To_X6Y12(ap_start_Boundary_X4Y12_To_X6Y12_out),
    .ap_rst_n_Boundary_X4Y12_To_X6Y12(ap_rst_n_Boundary_X4Y12_To_X6Y12_out),
    .ap_done_Boundary_X4Y12_To_X6Y12(ap_done_Boundary_X4Y12_To_X6Y12_in)
  );


  (* keep_hierarchy = "yes" *) CR_X6Y8_To_CR_X7Y9_ctrl CR_X6Y8_To_CR_X7Y9_ctrl_U0 (
    .PE_wrapper242_U0_fifo_w_out_V_V_din_pass_1(PE_wrapper242_U0_fifo_w_out_V_V_din_pass_1_in),
    .PE_wrapper242_U0_fifo_w_out_V_V_din_pass_2(PE_wrapper242_U0_fifo_w_out_V_V_din_pass_2_out),
    .fifo_w_PE_7_9_V_V_full_n_pass_1(fifo_w_PE_7_9_V_V_full_n_pass_1_out),
    .fifo_w_PE_7_9_V_V_full_n_pass_2(fifo_w_PE_7_9_V_V_full_n_pass_2_in),
    .PE_wrapper242_U0_fifo_w_out_V_V_write_pass_1(PE_wrapper242_U0_fifo_w_out_V_V_write_pass_1_in),
    .PE_wrapper242_U0_fifo_w_out_V_V_write_pass_2(PE_wrapper242_U0_fifo_w_out_V_V_write_pass_2_out),
    .cout_drain_IO_L1_out_wrapper474_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper474_U0_fifo_cout_drain_out_V_V_din_pass_0_in),
    .cout_drain_IO_L1_out_wrapper474_U0_fifo_cout_drain_out_V_V_din_pass_1(cout_drain_IO_L1_out_wrapper474_U0_fifo_cout_drain_out_V_V_din_pass_1_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_6_4_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_6_4_V_V_full_n_pass_0_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_6_4_V_V_full_n_pass_1(fifo_cout_drain_cout_drain_IO_L1_out_6_4_V_V_full_n_pass_1_in),
    .cout_drain_IO_L1_out_wrapper474_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper474_U0_fifo_cout_drain_out_V_V_write_pass_0_in),
    .cout_drain_IO_L1_out_wrapper474_U0_fifo_cout_drain_out_V_V_write_pass_1(cout_drain_IO_L1_out_wrapper474_U0_fifo_cout_drain_out_V_V_write_pass_1_out),
    .cout_drain_IO_L1_out_wrapper458_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper458_U0_fifo_cout_drain_out_V_V_din_pass_0_in),
    .cout_drain_IO_L1_out_wrapper458_U0_fifo_cout_drain_out_V_V_din_pass_1(cout_drain_IO_L1_out_wrapper458_U0_fifo_cout_drain_out_V_V_din_pass_1_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_5_4_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_5_4_V_V_full_n_pass_0_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_5_4_V_V_full_n_pass_1(fifo_cout_drain_cout_drain_IO_L1_out_5_4_V_V_full_n_pass_1_in),
    .cout_drain_IO_L1_out_wrapper458_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper458_U0_fifo_cout_drain_out_V_V_write_pass_0_in),
    .cout_drain_IO_L1_out_wrapper458_U0_fifo_cout_drain_out_V_V_write_pass_1(cout_drain_IO_L1_out_wrapper458_U0_fifo_cout_drain_out_V_V_write_pass_1_out),
    .PE_wrapper231_U0_fifo_cin_out_V_V_din_pass_3(PE_wrapper231_U0_fifo_cin_out_V_V_din_pass_3_in),
    .PE_wrapper231_U0_fifo_cin_out_V_V_din_pass_4(PE_wrapper231_U0_fifo_cin_out_V_V_din_pass_4_out),
    .fifo_cin_PE_7_9_V_V_full_n_pass_3(fifo_cin_PE_7_9_V_V_full_n_pass_3_out),
    .fifo_cin_PE_7_9_V_V_full_n_pass_4(fifo_cin_PE_7_9_V_V_full_n_pass_4_in),
    .PE_wrapper231_U0_fifo_cin_out_V_V_write_pass_3(PE_wrapper231_U0_fifo_cin_out_V_V_write_pass_3_in),
    .PE_wrapper231_U0_fifo_cin_out_V_V_write_pass_4(PE_wrapper231_U0_fifo_cin_out_V_V_write_pass_4_out),
    .PE_wrapper217_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper217_U0_fifo_w_out_V_V_din_pass_0_in),
    .PE_wrapper217_U0_fifo_w_out_V_V_din_pass_1(PE_wrapper217_U0_fifo_w_out_V_V_din_pass_1_out),
    .fifo_w_PE_5_8_V_V_full_n_pass_0(fifo_w_PE_5_8_V_V_full_n_pass_0_out),
    .fifo_w_PE_5_8_V_V_full_n_pass_1(fifo_w_PE_5_8_V_V_full_n_pass_1_in),
    .PE_wrapper217_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper217_U0_fifo_w_out_V_V_write_pass_0_in),
    .PE_wrapper217_U0_fifo_w_out_V_V_write_pass_1(PE_wrapper217_U0_fifo_w_out_V_V_write_pass_1_out),
    .PE_wrapper168_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper168_U0_fifo_w_out_V_V_din_pass_0_in),
    .fifo_w_PE_1_7_V_V_full_n_pass_0(fifo_w_PE_1_7_V_V_full_n_pass_0_out),
    .PE_wrapper168_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper168_U0_fifo_w_out_V_V_write_pass_0_in),
    .PE_wrapper193_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper193_U0_fifo_w_out_V_V_din_pass_0_out),
    .fifo_w_PE_3_8_V_V_full_n_pass_0(fifo_w_PE_3_8_V_V_full_n_pass_0_in),
    .PE_wrapper193_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper193_U0_fifo_w_out_V_V_write_pass_0_out),
    .PE_wrapper181_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper181_U0_fifo_w_out_V_V_din_pass_0_out),
    .fifo_w_PE_2_8_V_V_full_n_pass_0(fifo_w_PE_2_8_V_V_full_n_pass_0_in),
    .PE_wrapper181_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper181_U0_fifo_w_out_V_V_write_pass_0_out),
    .cout_drain_IO_L2_out561_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L2_out561_U0_fifo_cout_drain_out_V_V_din_pass_0_out),
    .fifo_cout_drain_cout_drain_IO_L2_out_7_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L2_out_7_V_V_full_n_pass_0_in),
    .cout_drain_IO_L2_out561_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L2_out561_U0_fifo_cout_drain_out_V_V_write_pass_0_out),
    .PE_wrapper169_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper169_U0_fifo_w_out_V_V_din_pass_0_out),
    .fifo_w_PE_1_8_V_V_full_n_pass_0(fifo_w_PE_1_8_V_V_full_n_pass_0_in),
    .PE_wrapper169_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper169_U0_fifo_w_out_V_V_write_pass_0_out),
    .cin_IO_L2_in130_U0_fifo_cin_out_V_V_din_pass_0(cin_IO_L2_in130_U0_fifo_cin_out_V_V_din_pass_0_in),
    .fifo_cin_cin_IO_L2_in_7_V_V_full_n_pass_0(fifo_cin_cin_IO_L2_in_7_V_V_full_n_pass_0_out),
    .cin_IO_L2_in130_U0_fifo_cin_out_V_V_write_pass_0(cin_IO_L2_in130_U0_fifo_cin_out_V_V_write_pass_0_in),
    .PE_wrapper205_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper205_U0_fifo_cin_out_V_V_din_pass_0_out),
    .fifo_cin_PE_5_7_V_V_full_n_pass_0(fifo_cin_PE_5_7_V_V_full_n_pass_0_in),
    .PE_wrapper205_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper205_U0_fifo_cin_out_V_V_write_pass_0_out),
    .cout_drain_IO_L1_out_wrapper490_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper490_U0_fifo_cout_drain_out_V_V_din_pass_0_in),
    .fifo_cout_drain_cout_drain_IO_L1_out_7_4_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_7_4_V_V_full_n_pass_0_out),
    .cout_drain_IO_L1_out_wrapper490_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper490_U0_fifo_cout_drain_out_V_V_write_pass_0_in),
    .cin_IO_L2_in131_U0_fifo_cin_out_V_V_din_pass_0(cin_IO_L2_in131_U0_fifo_cin_out_V_V_din_pass_0_out),
    .fifo_cin_cin_IO_L2_in_8_V_V_full_n_pass_0(fifo_cin_cin_IO_L2_in_8_V_V_full_n_pass_0_in),
    .cin_IO_L2_in131_U0_fifo_cin_out_V_V_write_pass_0(cin_IO_L2_in131_U0_fifo_cin_out_V_V_write_pass_0_out),
    .PE_wrapper156_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper156_U0_fifo_w_out_V_V_din_pass_0_in),
    .fifo_w_PE_0_7_V_V_full_n_pass_0(fifo_w_PE_0_7_V_V_full_n_pass_0_out),
    .PE_wrapper156_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper156_U0_fifo_w_out_V_V_write_pass_0_in),
    .PE_wrapper157_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper157_U0_fifo_w_out_V_V_din_pass_0_out),
    .fifo_w_PE_0_8_V_V_full_n_pass_0(fifo_w_PE_0_8_V_V_full_n_pass_0_in),
    .PE_wrapper157_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper157_U0_fifo_w_out_V_V_write_pass_0_out),
    .PE_wrapper192_U0_fifo_w_out_V_V_din_pass_1(PE_wrapper192_U0_fifo_w_out_V_V_din_pass_1_in),
    .fifo_w_PE_3_7_V_V_full_n_pass_1(fifo_w_PE_3_7_V_V_full_n_pass_1_out),
    .PE_wrapper192_U0_fifo_w_out_V_V_write_pass_1(PE_wrapper192_U0_fifo_w_out_V_V_write_pass_1_in),
    .cout_drain_IO_L2_out560_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L2_out560_U0_fifo_cout_drain_out_V_V_din_pass_0_in),
    .fifo_cout_drain_cout_drain_IO_L2_out_8_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L2_out_8_V_V_full_n_pass_0_out),
    .cout_drain_IO_L2_out560_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L2_out560_U0_fifo_cout_drain_out_V_V_write_pass_0_in),
    .cout_drain_IO_L3_out_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L3_out_U0_fifo_cout_drain_out_V_V_din_pass_0_out),
    .fifo_cout_drain_cout_drain_IO_L3_out_serialize_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L3_out_serialize_V_V_full_n_pass_0_in),
    .cout_drain_IO_L3_out_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L3_out_U0_fifo_cout_drain_out_V_V_write_pass_0_out),
    .PE_wrapper180_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper180_U0_fifo_w_out_V_V_din_pass_0_in),
    .fifo_w_PE_2_7_V_V_full_n_pass_0(fifo_w_PE_2_7_V_V_full_n_pass_0_out),
    .PE_wrapper180_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper180_U0_fifo_w_out_V_V_write_pass_0_in),
    .PE_wrapper205_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper205_U0_fifo_cout_drain_out_V_din_pass_0_out),
    .fifo_cout_drain_PE_4_7_V_full_n_pass_0(fifo_cout_drain_PE_4_7_V_full_n_pass_0_in),
    .PE_wrapper205_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper205_U0_fifo_cout_drain_out_V_write_pass_0_out),
    .PE_wrapper205_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper205_U0_fifo_w_out_V_V_din_pass_0_out),
    .fifo_w_PE_4_8_V_V_full_n_pass_0(fifo_w_PE_4_8_V_V_full_n_pass_0_in),
    .PE_wrapper205_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper205_U0_fifo_w_out_V_V_write_pass_0_out),
    .PE_wrapper204_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper204_U0_fifo_w_out_V_V_din_pass_0_in),
    .fifo_w_PE_4_7_V_V_full_n_pass_0(fifo_w_PE_4_7_V_V_full_n_pass_0_out),
    .PE_wrapper204_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper204_U0_fifo_w_out_V_V_write_pass_0_in),
    .cout_drain_IO_L2_out568_U0_fifo_cout_drain_out_V_V_din_pass_3(cout_drain_IO_L2_out568_U0_fifo_cout_drain_out_V_V_din_pass_3_in),
    .fifo_cout_drain_cout_drain_IO_L2_out_0_V_V_full_n_pass_3(fifo_cout_drain_cout_drain_IO_L2_out_0_V_V_full_n_pass_3_out),
    .cout_drain_IO_L2_out568_U0_fifo_cout_drain_out_V_V_write_pass_3(cout_drain_IO_L2_out568_U0_fifo_cout_drain_out_V_V_write_pass_3_in),
    .ap_clk(ap_clk),
    .ap_start_Boundary_X6Y8_To_X8Y8(ap_start_Boundary_X6Y8_To_X8Y8_in),
    .ap_rst_n_Boundary_X6Y8_To_X8Y8(ap_rst_n_Boundary_X6Y8_To_X8Y8_in),
    .ap_done_Boundary_X6Y8_To_X8Y8(ap_done_Boundary_X6Y8_To_X8Y8_out),
    .ap_start_Boundary_X6Y10_To_X8Y10(ap_start_Boundary_X6Y10_To_X8Y10_out),
    .ap_rst_n_Boundary_X6Y10_To_X8Y10(ap_rst_n_Boundary_X6Y10_To_X8Y10_out),
    .ap_done_Boundary_X6Y10_To_X8Y10(ap_done_Boundary_X6Y10_To_X8Y10_in)
  );


  (* keep_hierarchy = "yes" *) CR_X6Y10_To_CR_X7Y11_ctrl CR_X6Y10_To_CR_X7Y11_ctrl_U0 (
    .PE_wrapper242_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper242_U0_fifo_w_out_V_V_din_pass_0_in),
    .PE_wrapper242_U0_fifo_w_out_V_V_din_pass_1(PE_wrapper242_U0_fifo_w_out_V_V_din_pass_1_out),
    .fifo_w_PE_7_9_V_V_full_n_pass_0(fifo_w_PE_7_9_V_V_full_n_pass_0_out),
    .fifo_w_PE_7_9_V_V_full_n_pass_1(fifo_w_PE_7_9_V_V_full_n_pass_1_in),
    .PE_wrapper242_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper242_U0_fifo_w_out_V_V_write_pass_0_in),
    .PE_wrapper242_U0_fifo_w_out_V_V_write_pass_1(PE_wrapper242_U0_fifo_w_out_V_V_write_pass_1_out),
    .PE_wrapper231_U0_fifo_cin_out_V_V_din_pass_2(PE_wrapper231_U0_fifo_cin_out_V_V_din_pass_2_in),
    .PE_wrapper231_U0_fifo_cin_out_V_V_din_pass_3(PE_wrapper231_U0_fifo_cin_out_V_V_din_pass_3_out),
    .fifo_cin_PE_7_9_V_V_full_n_pass_2(fifo_cin_PE_7_9_V_V_full_n_pass_2_out),
    .fifo_cin_PE_7_9_V_V_full_n_pass_3(fifo_cin_PE_7_9_V_V_full_n_pass_3_in),
    .PE_wrapper231_U0_fifo_cin_out_V_V_write_pass_2(PE_wrapper231_U0_fifo_cin_out_V_V_write_pass_2_in),
    .PE_wrapper231_U0_fifo_cin_out_V_V_write_pass_3(PE_wrapper231_U0_fifo_cin_out_V_V_write_pass_3_out),
    .PE_wrapper158_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper158_U0_fifo_w_out_V_V_din_pass_0_out),
    .fifo_w_PE_0_9_V_V_full_n_pass_0(fifo_w_PE_0_9_V_V_full_n_pass_0_in),
    .PE_wrapper158_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper158_U0_fifo_w_out_V_V_write_pass_0_out),
    .PE_wrapper193_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper193_U0_fifo_w_out_V_V_din_pass_0_in),
    .fifo_w_PE_3_8_V_V_full_n_pass_0(fifo_w_PE_3_8_V_V_full_n_pass_0_out),
    .PE_wrapper193_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper193_U0_fifo_w_out_V_V_write_pass_0_in),
    .PE_wrapper170_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper170_U0_fifo_w_out_V_V_din_pass_0_out),
    .fifo_w_PE_1_9_V_V_full_n_pass_0(fifo_w_PE_1_9_V_V_full_n_pass_0_in),
    .PE_wrapper170_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper170_U0_fifo_w_out_V_V_write_pass_0_out),
    .cout_drain_IO_L2_out559_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L2_out559_U0_fifo_cout_drain_out_V_V_din_pass_0_in),
    .fifo_cout_drain_cout_drain_IO_L2_out_9_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L2_out_9_V_V_full_n_pass_0_out),
    .cout_drain_IO_L2_out559_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L2_out559_U0_fifo_cout_drain_out_V_V_write_pass_0_in),
    .PE_wrapper181_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper181_U0_fifo_w_out_V_V_din_pass_0_in),
    .fifo_w_PE_2_8_V_V_full_n_pass_0(fifo_w_PE_2_8_V_V_full_n_pass_0_out),
    .PE_wrapper181_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper181_U0_fifo_w_out_V_V_write_pass_0_in),
    .PE_wrapper206_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper206_U0_fifo_w_out_V_V_din_pass_0_out),
    .fifo_w_PE_4_9_V_V_full_n_pass_0(fifo_w_PE_4_9_V_V_full_n_pass_0_in),
    .PE_wrapper206_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper206_U0_fifo_w_out_V_V_write_pass_0_out),
    .cin_IO_L2_in132_U0_fifo_cin_out_V_V_din_pass_0(cin_IO_L2_in132_U0_fifo_cin_out_V_V_din_pass_0_out),
    .fifo_cin_cin_IO_L2_in_9_V_V_full_n_pass_0(fifo_cin_cin_IO_L2_in_9_V_V_full_n_pass_0_in),
    .cin_IO_L2_in132_U0_fifo_cin_out_V_V_write_pass_0(cin_IO_L2_in132_U0_fifo_cin_out_V_V_write_pass_0_out),
    .PE_wrapper218_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper218_U0_fifo_cout_drain_out_V_din_pass_0_out),
    .fifo_cout_drain_PE_5_8_V_full_n_pass_0(fifo_cout_drain_PE_5_8_V_full_n_pass_0_in),
    .PE_wrapper218_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper218_U0_fifo_cout_drain_out_V_write_pass_0_out),
    .cout_drain_IO_L1_out_wrapper506_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper506_U0_fifo_cout_drain_out_V_V_din_pass_0_in),
    .fifo_cout_drain_cout_drain_IO_L1_out_8_4_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_8_4_V_V_full_n_pass_0_out),
    .cout_drain_IO_L1_out_wrapper506_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper506_U0_fifo_cout_drain_out_V_V_write_pass_0_in),
    .PE_wrapper169_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper169_U0_fifo_w_out_V_V_din_pass_0_in),
    .fifo_w_PE_1_8_V_V_full_n_pass_0(fifo_w_PE_1_8_V_V_full_n_pass_0_out),
    .PE_wrapper169_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper169_U0_fifo_w_out_V_V_write_pass_0_in),
    .PE_wrapper217_U0_fifo_w_out_V_V_din_pass_1(PE_wrapper217_U0_fifo_w_out_V_V_din_pass_1_in),
    .fifo_w_PE_5_8_V_V_full_n_pass_1(fifo_w_PE_5_8_V_V_full_n_pass_1_out),
    .PE_wrapper217_U0_fifo_w_out_V_V_write_pass_1(PE_wrapper217_U0_fifo_w_out_V_V_write_pass_1_in),
    .cin_IO_L2_in131_U0_fifo_cin_out_V_V_din_pass_0(cin_IO_L2_in131_U0_fifo_cin_out_V_V_din_pass_0_in),
    .fifo_cin_cin_IO_L2_in_8_V_V_full_n_pass_0(fifo_cin_cin_IO_L2_in_8_V_V_full_n_pass_0_out),
    .cin_IO_L2_in131_U0_fifo_cin_out_V_V_write_pass_0(cin_IO_L2_in131_U0_fifo_cin_out_V_V_write_pass_0_in),
    .PE_wrapper157_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper157_U0_fifo_w_out_V_V_din_pass_0_in),
    .fifo_w_PE_0_8_V_V_full_n_pass_0(fifo_w_PE_0_8_V_V_full_n_pass_0_out),
    .PE_wrapper157_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper157_U0_fifo_w_out_V_V_write_pass_0_in),
    .PE_wrapper182_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper182_U0_fifo_w_out_V_V_din_pass_0_out),
    .fifo_w_PE_2_9_V_V_full_n_pass_0(fifo_w_PE_2_9_V_V_full_n_pass_0_in),
    .PE_wrapper182_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper182_U0_fifo_w_out_V_V_write_pass_0_out),
    .cout_drain_IO_L2_out560_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L2_out560_U0_fifo_cout_drain_out_V_V_din_pass_0_out),
    .fifo_cout_drain_cout_drain_IO_L2_out_8_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L2_out_8_V_V_full_n_pass_0_in),
    .cout_drain_IO_L2_out560_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L2_out560_U0_fifo_cout_drain_out_V_V_write_pass_0_out),
    .PE_wrapper205_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper205_U0_fifo_w_out_V_V_din_pass_0_in),
    .fifo_w_PE_4_8_V_V_full_n_pass_0(fifo_w_PE_4_8_V_V_full_n_pass_0_out),
    .PE_wrapper205_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper205_U0_fifo_w_out_V_V_write_pass_0_in),
    .PE_wrapper218_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper218_U0_fifo_w_out_V_V_din_pass_0_out),
    .fifo_w_PE_5_9_V_V_full_n_pass_0(fifo_w_PE_5_9_V_V_full_n_pass_0_in),
    .PE_wrapper218_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper218_U0_fifo_w_out_V_V_write_pass_0_out),
    .PE_wrapper206_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper206_U0_fifo_cout_drain_out_V_din_pass_0_out),
    .fifo_cout_drain_PE_4_8_V_full_n_pass_0(fifo_cout_drain_PE_4_8_V_full_n_pass_0_in),
    .PE_wrapper206_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper206_U0_fifo_cout_drain_out_V_write_pass_0_out),
    .PE_wrapper218_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper218_U0_fifo_cin_out_V_V_din_pass_0_out),
    .fifo_cin_PE_6_8_V_V_full_n_pass_0(fifo_cin_PE_6_8_V_V_full_n_pass_0_in),
    .PE_wrapper218_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper218_U0_fifo_cin_out_V_V_write_pass_0_out),
    .PE_wrapper194_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper194_U0_fifo_w_out_V_V_din_pass_0_out),
    .fifo_w_PE_3_9_V_V_full_n_pass_0(fifo_w_PE_3_9_V_V_full_n_pass_0_in),
    .PE_wrapper194_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper194_U0_fifo_w_out_V_V_write_pass_0_out),
    .ap_clk(ap_clk),
    .ap_start_Boundary_X6Y10_To_X8Y10(ap_start_Boundary_X6Y10_To_X8Y10_in),
    .ap_rst_n_Boundary_X6Y10_To_X8Y10(ap_rst_n_Boundary_X6Y10_To_X8Y10_in),
    .ap_done_Boundary_X6Y10_To_X8Y10(ap_done_Boundary_X6Y10_To_X8Y10_out),
    .ap_start_Boundary_X6Y12_To_X8Y12(ap_start_Boundary_X6Y12_To_X8Y12_out),
    .ap_rst_n_Boundary_X6Y12_To_X8Y12(ap_rst_n_Boundary_X6Y12_To_X8Y12_out),
    .ap_done_Boundary_X6Y12_To_X8Y12(ap_done_Boundary_X6Y12_To_X8Y12_in)
  );


  (* keep_hierarchy = "yes" *) CR_X4Y14_To_CR_X5Y15_ctrl CR_X4Y14_To_CR_X5Y15_ctrl_U0 (
    .PE_wrapper256_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper256_U0_fifo_cin_out_V_V_din_pass_0_in),
    .PE_wrapper256_U0_fifo_cin_out_V_V_din_pass_1(PE_wrapper256_U0_fifo_cin_out_V_V_din_pass_1_out),
    .fifo_cin_PE_9_10_V_V_full_n_pass_0(fifo_cin_PE_9_10_V_V_full_n_pass_0_out),
    .fifo_cin_PE_9_10_V_V_full_n_pass_1(fifo_cin_PE_9_10_V_V_full_n_pass_1_in),
    .PE_wrapper256_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper256_U0_fifo_cin_out_V_V_write_pass_0_in),
    .PE_wrapper256_U0_fifo_cin_out_V_V_write_pass_1(PE_wrapper256_U0_fifo_cin_out_V_V_write_pass_1_out),
    .PE_wrapper257_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper257_U0_fifo_cin_out_V_V_din_pass_0_in),
    .PE_wrapper257_U0_fifo_cin_out_V_V_din_pass_1(PE_wrapper257_U0_fifo_cin_out_V_V_din_pass_1_out),
    .fifo_cin_PE_9_11_V_V_full_n_pass_0(fifo_cin_PE_9_11_V_V_full_n_pass_0_out),
    .fifo_cin_PE_9_11_V_V_full_n_pass_1(fifo_cin_PE_9_11_V_V_full_n_pass_1_in),
    .PE_wrapper257_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper257_U0_fifo_cin_out_V_V_write_pass_0_in),
    .PE_wrapper257_U0_fifo_cin_out_V_V_write_pass_1(PE_wrapper257_U0_fifo_cin_out_V_V_write_pass_1_out),
    .cout_drain_IO_L1_out_wrapper551_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper551_U0_fifo_cout_drain_out_V_V_din_pass_0_in),
    .cout_drain_IO_L1_out_wrapper551_U0_fifo_cout_drain_out_V_V_din_pass_1(cout_drain_IO_L1_out_wrapper551_U0_fifo_cout_drain_out_V_V_din_pass_1_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_11_6_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_11_6_V_V_full_n_pass_0_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_11_6_V_V_full_n_pass_1(fifo_cout_drain_cout_drain_IO_L1_out_11_6_V_V_full_n_pass_1_in),
    .cout_drain_IO_L1_out_wrapper551_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper551_U0_fifo_cout_drain_out_V_V_write_pass_0_in),
    .cout_drain_IO_L1_out_wrapper551_U0_fifo_cout_drain_out_V_V_write_pass_1(cout_drain_IO_L1_out_wrapper551_U0_fifo_cout_drain_out_V_V_write_pass_1_out),
    .PE_wrapper161_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper161_U0_fifo_cin_out_V_V_din_pass_0_in),
    .PE_wrapper161_U0_fifo_cin_out_V_V_din_pass_1(PE_wrapper161_U0_fifo_cin_out_V_V_din_pass_1_out),
    .fifo_cin_PE_1_11_V_V_full_n_pass_0(fifo_cin_PE_1_11_V_V_full_n_pass_0_out),
    .fifo_cin_PE_1_11_V_V_full_n_pass_1(fifo_cin_PE_1_11_V_V_full_n_pass_1_in),
    .PE_wrapper161_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper161_U0_fifo_cin_out_V_V_write_pass_0_in),
    .PE_wrapper161_U0_fifo_cin_out_V_V_write_pass_1(PE_wrapper161_U0_fifo_cin_out_V_V_write_pass_1_out),
    .PE_wrapper185_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper185_U0_fifo_cout_drain_out_V_din_pass_0_in),
    .PE_wrapper185_U0_fifo_cout_drain_out_V_din_pass_1(PE_wrapper185_U0_fifo_cout_drain_out_V_din_pass_1_out),
    .fifo_cout_drain_PE_2_11_V_full_n_pass_0(fifo_cout_drain_PE_2_11_V_full_n_pass_0_out),
    .fifo_cout_drain_PE_2_11_V_full_n_pass_1(fifo_cout_drain_PE_2_11_V_full_n_pass_1_in),
    .PE_wrapper185_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper185_U0_fifo_cout_drain_out_V_write_pass_0_in),
    .PE_wrapper185_U0_fifo_cout_drain_out_V_write_pass_1(PE_wrapper185_U0_fifo_cout_drain_out_V_write_pass_1_out),
    .cout_drain_IO_L1_out_wrapper518_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper518_U0_fifo_cout_drain_out_V_V_din_pass_0_in),
    .cout_drain_IO_L1_out_wrapper518_U0_fifo_cout_drain_out_V_V_din_pass_1(cout_drain_IO_L1_out_wrapper518_U0_fifo_cout_drain_out_V_V_din_pass_1_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_9_8_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_9_8_V_V_full_n_pass_0_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_9_8_V_V_full_n_pass_1(fifo_cout_drain_cout_drain_IO_L1_out_9_8_V_V_full_n_pass_1_in),
    .cout_drain_IO_L1_out_wrapper518_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper518_U0_fifo_cout_drain_out_V_V_write_pass_0_in),
    .cout_drain_IO_L1_out_wrapper518_U0_fifo_cout_drain_out_V_V_write_pass_1(cout_drain_IO_L1_out_wrapper518_U0_fifo_cout_drain_out_V_V_write_pass_1_out),
    .cout_drain_IO_L1_out_wrapper534_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper534_U0_fifo_cout_drain_out_V_V_din_pass_0_in),
    .cout_drain_IO_L1_out_wrapper534_U0_fifo_cout_drain_out_V_V_din_pass_1(cout_drain_IO_L1_out_wrapper534_U0_fifo_cout_drain_out_V_V_din_pass_1_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_10_8_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_10_8_V_V_full_n_pass_0_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_10_8_V_V_full_n_pass_1(fifo_cout_drain_cout_drain_IO_L1_out_10_8_V_V_full_n_pass_1_in),
    .cout_drain_IO_L1_out_wrapper534_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper534_U0_fifo_cout_drain_out_V_V_write_pass_0_in),
    .cout_drain_IO_L1_out_wrapper534_U0_fifo_cout_drain_out_V_V_write_pass_1(cout_drain_IO_L1_out_wrapper534_U0_fifo_cout_drain_out_V_V_write_pass_1_out),
    .PE_wrapper197_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper197_U0_fifo_cout_drain_out_V_din_pass_0_in),
    .PE_wrapper197_U0_fifo_cout_drain_out_V_din_pass_1(PE_wrapper197_U0_fifo_cout_drain_out_V_din_pass_1_out),
    .fifo_cout_drain_PE_3_11_V_full_n_pass_0(fifo_cout_drain_PE_3_11_V_full_n_pass_0_out),
    .fifo_cout_drain_PE_3_11_V_full_n_pass_1(fifo_cout_drain_PE_3_11_V_full_n_pass_1_in),
    .PE_wrapper197_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper197_U0_fifo_cout_drain_out_V_write_pass_0_in),
    .PE_wrapper197_U0_fifo_cout_drain_out_V_write_pass_1(PE_wrapper197_U0_fifo_cout_drain_out_V_write_pass_1_out),
    .cout_drain_IO_L1_out_wrapper523_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper523_U0_fifo_cout_drain_out_V_V_din_pass_0_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_9_3_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_9_3_V_V_full_n_pass_0_in),
    .cout_drain_IO_L1_out_wrapper523_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper523_U0_fifo_cout_drain_out_V_V_write_pass_0_out),
    .cout_drain_IO_L1_out_wrapper535_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper535_U0_fifo_cout_drain_out_V_V_din_pass_0_in),
    .fifo_cout_drain_cout_drain_IO_L1_out_10_7_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_10_7_V_V_full_n_pass_0_out),
    .cout_drain_IO_L1_out_wrapper535_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper535_U0_fifo_cout_drain_out_V_V_write_pass_0_in),
    .cout_drain_IO_L1_out_wrapper537_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper537_U0_fifo_cout_drain_out_V_V_din_pass_0_in),
    .fifo_cout_drain_cout_drain_IO_L1_out_10_5_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_10_5_V_V_full_n_pass_0_out),
    .cout_drain_IO_L1_out_wrapper537_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper537_U0_fifo_cout_drain_out_V_V_write_pass_0_in),
    .cout_drain_IO_L1_out_wrapper555_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper555_U0_fifo_cout_drain_out_V_V_din_pass_0_in),
    .fifo_cout_drain_cout_drain_IO_L1_out_11_2_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_11_2_V_V_full_n_pass_0_out),
    .cout_drain_IO_L1_out_wrapper555_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper555_U0_fifo_cout_drain_out_V_V_write_pass_0_in),
    .PE_wrapper196_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper196_U0_fifo_cin_out_V_V_din_pass_0_out),
    .fifo_cin_PE_4_10_V_V_full_n_pass_0(fifo_cin_PE_4_10_V_V_full_n_pass_0_in),
    .PE_wrapper196_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper196_U0_fifo_cin_out_V_V_write_pass_0_out),
    .cout_drain_IO_L1_out_wrapper556_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper556_U0_fifo_cout_drain_out_V_V_din_pass_0_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_11_1_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_11_1_V_V_full_n_pass_0_in),
    .cout_drain_IO_L1_out_wrapper556_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper556_U0_fifo_cout_drain_out_V_V_write_pass_0_out),
    .cout_drain_IO_L1_out_wrapper539_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper539_U0_fifo_cout_drain_out_V_V_din_pass_0_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_10_3_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_10_3_V_V_full_n_pass_0_in),
    .cout_drain_IO_L1_out_wrapper539_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper539_U0_fifo_cout_drain_out_V_V_write_pass_0_out),
    .PE_wrapper231_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper231_U0_fifo_w_out_V_V_din_pass_0_out),
    .fifo_w_PE_6_10_V_V_full_n_pass_0(fifo_w_PE_6_10_V_V_full_n_pass_0_in),
    .PE_wrapper231_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper231_U0_fifo_w_out_V_V_write_pass_0_out),
    .PE_wrapper231_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper231_U0_fifo_cout_drain_out_V_din_pass_0_out),
    .fifo_cout_drain_PE_6_9_V_full_n_pass_0(fifo_cout_drain_PE_6_9_V_full_n_pass_0_in),
    .PE_wrapper231_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper231_U0_fifo_cout_drain_out_V_write_pass_0_out),
    .PE_wrapper230_U0_fifo_w_out_V_V_din_pass_1(PE_wrapper230_U0_fifo_w_out_V_V_din_pass_1_in),
    .fifo_w_PE_6_9_V_V_full_n_pass_1(fifo_w_PE_6_9_V_V_full_n_pass_1_out),
    .PE_wrapper230_U0_fifo_w_out_V_V_write_pass_1(PE_wrapper230_U0_fifo_w_out_V_V_write_pass_1_in),
    .cout_drain_IO_L2_out558_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L2_out558_U0_fifo_cout_drain_out_V_V_din_pass_0_out),
    .fifo_cout_drain_cout_drain_IO_L2_out_10_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L2_out_10_V_V_full_n_pass_0_in),
    .cout_drain_IO_L2_out558_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L2_out558_U0_fifo_cout_drain_out_V_V_write_pass_0_out),
    .PE_wrapper221_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper221_U0_fifo_cout_drain_out_V_din_pass_0_out),
    .fifo_cout_drain_PE_5_11_V_full_n_pass_0(fifo_cout_drain_PE_5_11_V_full_n_pass_0_in),
    .PE_wrapper221_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper221_U0_fifo_cout_drain_out_V_write_pass_0_out),
    .PE_wrapper184_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper184_U0_fifo_w_out_V_V_din_pass_0_out),
    .fifo_w_PE_2_11_V_V_full_n_pass_0(fifo_w_PE_2_11_V_V_full_n_pass_0_in),
    .PE_wrapper184_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper184_U0_fifo_w_out_V_V_write_pass_0_out),
    .PE_wrapper232_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper232_U0_fifo_cout_drain_out_V_din_pass_0_in),
    .fifo_cout_drain_PE_6_10_V_full_n_pass_0(fifo_cout_drain_PE_6_10_V_full_n_pass_0_out),
    .PE_wrapper232_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper232_U0_fifo_cout_drain_out_V_write_pass_0_in),
    .cout_drain_IO_L1_out_wrapper522_U0_fifo_cout_drain_out_V_V_din_pass_1(cout_drain_IO_L1_out_wrapper522_U0_fifo_cout_drain_out_V_V_din_pass_1_in),
    .fifo_cout_drain_cout_drain_IO_L1_out_9_4_V_V_full_n_pass_1(fifo_cout_drain_cout_drain_IO_L1_out_9_4_V_V_full_n_pass_1_out),
    .cout_drain_IO_L1_out_wrapper522_U0_fifo_cout_drain_out_V_V_write_pass_1(cout_drain_IO_L1_out_wrapper522_U0_fifo_cout_drain_out_V_V_write_pass_1_in),
    .PE_wrapper196_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper196_U0_fifo_w_out_V_V_din_pass_0_out),
    .fifo_w_PE_3_11_V_V_full_n_pass_0(fifo_w_PE_3_11_V_V_full_n_pass_0_in),
    .PE_wrapper196_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper196_U0_fifo_w_out_V_V_write_pass_0_out),
    .PE_wrapper209_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper209_U0_fifo_w_out_V_V_din_pass_0_out),
    .fifo_w_PE_4_12_V_V_full_n_pass_0(fifo_w_PE_4_12_V_V_full_n_pass_0_in),
    .PE_wrapper209_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper209_U0_fifo_w_out_V_V_write_pass_0_out),
    .cout_drain_IO_L1_out_wrapper552_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper552_U0_fifo_cout_drain_out_V_V_din_pass_0_in),
    .fifo_cout_drain_cout_drain_IO_L1_out_11_5_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_11_5_V_V_full_n_pass_0_out),
    .cout_drain_IO_L1_out_wrapper552_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper552_U0_fifo_cout_drain_out_V_V_write_pass_0_in),
    .PE_wrapper233_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper233_U0_fifo_cin_out_V_V_din_pass_0_out),
    .fifo_cin_PE_7_11_V_V_full_n_pass_0(fifo_cin_PE_7_11_V_V_full_n_pass_0_in),
    .PE_wrapper233_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper233_U0_fifo_cin_out_V_V_write_pass_0_out),
    .PE_wrapper184_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper184_U0_fifo_cout_drain_out_V_din_pass_0_out),
    .fifo_cout_drain_PE_2_10_V_full_n_pass_0(fifo_cout_drain_PE_2_10_V_full_n_pass_0_in),
    .PE_wrapper184_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper184_U0_fifo_cout_drain_out_V_write_pass_0_out),
    .cout_drain_IO_L2_out_boundary_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L2_out_boundary_U0_fifo_cout_drain_out_V_V_din_pass_0_in),
    .fifo_cout_drain_cout_drain_IO_L2_out_11_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L2_out_11_V_V_full_n_pass_0_out),
    .cout_drain_IO_L2_out_boundary_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L2_out_boundary_U0_fifo_cout_drain_out_V_V_write_pass_0_in),
    .PE_wrapper197_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper197_U0_fifo_cin_out_V_V_din_pass_0_in),
    .fifo_cin_PE_4_11_V_V_full_n_pass_0(fifo_cin_PE_4_11_V_V_full_n_pass_0_out),
    .PE_wrapper197_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper197_U0_fifo_cin_out_V_V_write_pass_0_in),
    .cout_drain_IO_L1_out_wrapper542_U0_fifo_cout_drain_out_V_V_din_pass_1(cout_drain_IO_L1_out_wrapper542_U0_fifo_cout_drain_out_V_V_din_pass_1_in),
    .fifo_cout_drain_cout_drain_IO_L1_out_10_0_V_V_full_n_pass_1(fifo_cout_drain_cout_drain_IO_L1_out_10_0_V_V_full_n_pass_1_out),
    .cout_drain_IO_L1_out_wrapper542_U0_fifo_cout_drain_out_V_V_write_pass_1(cout_drain_IO_L1_out_wrapper542_U0_fifo_cout_drain_out_V_V_write_pass_1_in),
    .PE_wrapper219_U0_fifo_cin_out_V_V_din_pass_1(PE_wrapper219_U0_fifo_cin_out_V_V_din_pass_1_in),
    .fifo_cin_PE_6_9_V_V_full_n_pass_1(fifo_cin_PE_6_9_V_V_full_n_pass_1_out),
    .PE_wrapper219_U0_fifo_cin_out_V_V_write_pass_1(PE_wrapper219_U0_fifo_cin_out_V_V_write_pass_1_in),
    .PE_wrapper173_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper173_U0_fifo_cout_drain_out_V_din_pass_0_in),
    .fifo_cout_drain_PE_1_11_V_full_n_pass_0(fifo_cout_drain_PE_1_11_V_full_n_pass_0_out),
    .PE_wrapper173_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper173_U0_fifo_cout_drain_out_V_write_pass_0_in),
    .cout_drain_IO_L1_out_wrapper549_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper549_U0_fifo_cout_drain_out_V_V_din_pass_0_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_11_8_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_11_8_V_V_full_n_pass_0_in),
    .cout_drain_IO_L1_out_wrapper549_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper549_U0_fifo_cout_drain_out_V_V_write_pass_0_out),
    .PE_wrapper172_U0_fifo_cin_out_V_V_din_pass_1(PE_wrapper172_U0_fifo_cin_out_V_V_din_pass_1_in),
    .fifo_cin_PE_2_10_V_V_full_n_pass_1(fifo_cin_PE_2_10_V_V_full_n_pass_1_out),
    .PE_wrapper172_U0_fifo_cin_out_V_V_write_pass_1(PE_wrapper172_U0_fifo_cin_out_V_V_write_pass_1_in),
    .PE_wrapper195_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper195_U0_fifo_cin_out_V_V_din_pass_0_out),
    .fifo_cin_PE_4_9_V_V_full_n_pass_0(fifo_cin_PE_4_9_V_V_full_n_pass_0_in),
    .PE_wrapper195_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper195_U0_fifo_cin_out_V_V_write_pass_0_out),
    .cout_drain_IO_L1_out_wrapper536_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper536_U0_fifo_cout_drain_out_V_V_din_pass_0_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_10_6_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_10_6_V_V_full_n_pass_0_in),
    .cout_drain_IO_L1_out_wrapper536_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper536_U0_fifo_cout_drain_out_V_V_write_pass_0_out),
    .PE_wrapper208_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper208_U0_fifo_cout_drain_out_V_din_pass_0_in),
    .fifo_cout_drain_PE_4_10_V_full_n_pass_0(fifo_cout_drain_PE_4_10_V_full_n_pass_0_out),
    .PE_wrapper208_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper208_U0_fifo_cout_drain_out_V_write_pass_0_in),
    .PE_wrapper220_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper220_U0_fifo_w_out_V_V_din_pass_0_in),
    .fifo_w_PE_5_11_V_V_full_n_pass_0(fifo_w_PE_5_11_V_V_full_n_pass_0_out),
    .PE_wrapper220_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper220_U0_fifo_w_out_V_V_write_pass_0_in),
    .cin_IO_L2_in134_U0_fifo_cin_out_V_V_din_pass_1(cin_IO_L2_in134_U0_fifo_cin_out_V_V_din_pass_1_in),
    .fifo_cin_cin_IO_L2_in_11_V_V_full_n_pass_1(fifo_cin_cin_IO_L2_in_11_V_V_full_n_pass_1_out),
    .cin_IO_L2_in134_U0_fifo_cin_out_V_V_write_pass_1(cin_IO_L2_in134_U0_fifo_cin_out_V_V_write_pass_1_in),
    .cout_drain_IO_L1_out_wrapper520_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper520_U0_fifo_cout_drain_out_V_V_din_pass_0_in),
    .fifo_cout_drain_cout_drain_IO_L1_out_9_6_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_9_6_V_V_full_n_pass_0_out),
    .cout_drain_IO_L1_out_wrapper520_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper520_U0_fifo_cout_drain_out_V_V_write_pass_0_in),
    .PE_wrapper257_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper257_U0_fifo_cout_drain_out_V_din_pass_0_in),
    .fifo_cout_drain_PE_8_11_V_full_n_pass_0(fifo_cout_drain_PE_8_11_V_full_n_pass_0_out),
    .PE_wrapper257_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper257_U0_fifo_cout_drain_out_V_write_pass_0_in),
    .cin_IO_L2_in_boundary_U0_fifo_cin_local_out_V_V_din_pass_0(cin_IO_L2_in_boundary_U0_fifo_cin_local_out_V_V_din_pass_0_out),
    .fifo_cin_PE_0_11_V_V_full_n_pass_0(fifo_cin_PE_0_11_V_V_full_n_pass_0_in),
    .cin_IO_L2_in_boundary_U0_fifo_cin_local_out_V_V_write_pass_0(cin_IO_L2_in_boundary_U0_fifo_cin_local_out_V_V_write_pass_0_out),
    .PE_wrapper232_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper232_U0_fifo_w_out_V_V_din_pass_0_in),
    .fifo_w_PE_6_11_V_V_full_n_pass_0(fifo_w_PE_6_11_V_V_full_n_pass_0_out),
    .PE_wrapper232_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper232_U0_fifo_w_out_V_V_write_pass_0_in),
    .PE_wrapper183_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper183_U0_fifo_w_out_V_V_din_pass_0_in),
    .fifo_w_PE_2_10_V_V_full_n_pass_0(fifo_w_PE_2_10_V_V_full_n_pass_0_out),
    .PE_wrapper183_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper183_U0_fifo_w_out_V_V_write_pass_0_in),
    .PE_wrapper221_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper221_U0_fifo_w_out_V_V_din_pass_0_out),
    .fifo_w_PE_5_12_V_V_full_n_pass_0(fifo_w_PE_5_12_V_V_full_n_pass_0_in),
    .PE_wrapper221_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper221_U0_fifo_w_out_V_V_write_pass_0_out),
    .PE_wrapper208_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper208_U0_fifo_w_out_V_V_din_pass_0_in),
    .fifo_w_PE_4_11_V_V_full_n_pass_0(fifo_w_PE_4_11_V_V_full_n_pass_0_out),
    .PE_wrapper208_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper208_U0_fifo_w_out_V_V_write_pass_0_in),
    .PE_wrapper233_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper233_U0_fifo_cout_drain_out_V_din_pass_0_out),
    .fifo_cout_drain_PE_6_11_V_full_n_pass_0(fifo_cout_drain_PE_6_11_V_full_n_pass_0_in),
    .PE_wrapper233_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper233_U0_fifo_cout_drain_out_V_write_pass_0_out),
    .PE_wrapper183_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper183_U0_fifo_cin_out_V_V_din_pass_0_in),
    .fifo_cin_PE_3_9_V_V_full_n_pass_0(fifo_cin_PE_3_9_V_V_full_n_pass_0_out),
    .PE_wrapper183_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper183_U0_fifo_cin_out_V_V_write_pass_0_in),
    .PE_wrapper194_U0_fifo_w_out_V_V_din_pass_2(PE_wrapper194_U0_fifo_w_out_V_V_din_pass_2_in),
    .fifo_w_PE_3_9_V_V_full_n_pass_2(fifo_w_PE_3_9_V_V_full_n_pass_2_out),
    .PE_wrapper194_U0_fifo_w_out_V_V_write_pass_2(PE_wrapper194_U0_fifo_w_out_V_V_write_pass_2_in),
    .PE_wrapper231_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper231_U0_fifo_cin_out_V_V_din_pass_0_out),
    .fifo_cin_PE_7_9_V_V_full_n_pass_0(fifo_cin_PE_7_9_V_V_full_n_pass_0_in),
    .PE_wrapper231_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper231_U0_fifo_cin_out_V_V_write_pass_0_out),
    .PE_wrapper185_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper185_U0_fifo_w_out_V_V_din_pass_0_in),
    .fifo_w_PE_2_12_V_V_full_n_pass_0(fifo_w_PE_2_12_V_V_full_n_pass_0_out),
    .PE_wrapper185_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper185_U0_fifo_w_out_V_V_write_pass_0_in),
    .cout_drain_IO_L1_out_wrapper548_U0_fifo_cout_drain_out_V_V_din_pass_1(cout_drain_IO_L1_out_wrapper548_U0_fifo_cout_drain_out_V_V_din_pass_1_in),
    .fifo_cout_drain_cout_drain_IO_L1_out_11_9_V_V_full_n_pass_1(fifo_cout_drain_cout_drain_IO_L1_out_11_9_V_V_full_n_pass_1_out),
    .cout_drain_IO_L1_out_wrapper548_U0_fifo_cout_drain_out_V_V_write_pass_1(cout_drain_IO_L1_out_wrapper548_U0_fifo_cout_drain_out_V_V_write_pass_1_in),
    .cout_drain_IO_L1_out_wrapper521_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper521_U0_fifo_cout_drain_out_V_V_din_pass_0_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_9_5_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_9_5_V_V_full_n_pass_0_in),
    .cout_drain_IO_L1_out_wrapper521_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper521_U0_fifo_cout_drain_out_V_V_write_pass_0_out),
    .PE_wrapper219_U0_fifo_cout_drain_out_V_din_pass_1(PE_wrapper219_U0_fifo_cout_drain_out_V_din_pass_1_in),
    .fifo_cout_drain_PE_5_9_V_full_n_pass_1(fifo_cout_drain_PE_5_9_V_full_n_pass_1_out),
    .PE_wrapper219_U0_fifo_cout_drain_out_V_write_pass_1(PE_wrapper219_U0_fifo_cout_drain_out_V_write_pass_1_in),
    .cout_drain_IO_L1_out_wrapper553_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper553_U0_fifo_cout_drain_out_V_V_din_pass_0_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_11_4_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_11_4_V_V_full_n_pass_0_in),
    .cout_drain_IO_L1_out_wrapper553_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper553_U0_fifo_cout_drain_out_V_V_write_pass_0_out),
    .ap_clk(ap_clk),
    .ap_start_Boundary_X4Y14_To_X6Y14(ap_start_Boundary_X4Y14_To_X6Y14_in),
    .ap_rst_n_Boundary_X4Y14_To_X6Y14(ap_rst_n_Boundary_X4Y14_To_X6Y14_in),
    .ap_done_Boundary_X4Y14_To_X6Y14(ap_done_Boundary_X4Y14_To_X6Y14_out)
  );


  (* keep_hierarchy = "yes" *) CR_X6Y12_To_CR_X7Y13_ctrl CR_X6Y12_To_CR_X7Y13_ctrl_U0 (
    .PE_wrapper231_U0_fifo_cin_out_V_V_din_pass_1(PE_wrapper231_U0_fifo_cin_out_V_V_din_pass_1_in),
    .PE_wrapper231_U0_fifo_cin_out_V_V_din_pass_2(PE_wrapper231_U0_fifo_cin_out_V_V_din_pass_2_out),
    .fifo_cin_PE_7_9_V_V_full_n_pass_1(fifo_cin_PE_7_9_V_V_full_n_pass_1_out),
    .fifo_cin_PE_7_9_V_V_full_n_pass_2(fifo_cin_PE_7_9_V_V_full_n_pass_2_in),
    .PE_wrapper231_U0_fifo_cin_out_V_V_write_pass_1(PE_wrapper231_U0_fifo_cin_out_V_V_write_pass_1_in),
    .PE_wrapper231_U0_fifo_cin_out_V_V_write_pass_2(PE_wrapper231_U0_fifo_cin_out_V_V_write_pass_2_out),
    .PE_wrapper244_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper244_U0_fifo_cin_out_V_V_din_pass_0_in),
    .PE_wrapper244_U0_fifo_cin_out_V_V_din_pass_1(PE_wrapper244_U0_fifo_cin_out_V_V_din_pass_1_out),
    .fifo_cin_PE_8_10_V_V_full_n_pass_0(fifo_cin_PE_8_10_V_V_full_n_pass_0_out),
    .fifo_cin_PE_8_10_V_V_full_n_pass_1(fifo_cin_PE_8_10_V_V_full_n_pass_1_in),
    .PE_wrapper244_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper244_U0_fifo_cin_out_V_V_write_pass_0_in),
    .PE_wrapper244_U0_fifo_cin_out_V_V_write_pass_1(PE_wrapper244_U0_fifo_cin_out_V_V_write_pass_1_out),
    .PE_wrapper173_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper173_U0_fifo_w_out_V_V_din_pass_0_in),
    .PE_wrapper173_U0_fifo_w_out_V_V_din_pass_1(PE_wrapper173_U0_fifo_w_out_V_V_din_pass_1_out),
    .fifo_w_PE_1_12_V_V_full_n_pass_0(fifo_w_PE_1_12_V_V_full_n_pass_0_out),
    .fifo_w_PE_1_12_V_V_full_n_pass_1(fifo_w_PE_1_12_V_V_full_n_pass_1_in),
    .PE_wrapper173_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper173_U0_fifo_w_out_V_V_write_pass_0_in),
    .PE_wrapper173_U0_fifo_w_out_V_V_write_pass_1(PE_wrapper173_U0_fifo_w_out_V_V_write_pass_1_out),
    .PE_wrapper255_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper255_U0_fifo_cout_drain_out_V_din_pass_0_in),
    .PE_wrapper255_U0_fifo_cout_drain_out_V_din_pass_1(PE_wrapper255_U0_fifo_cout_drain_out_V_din_pass_1_out),
    .fifo_cout_drain_PE_8_9_V_full_n_pass_0(fifo_cout_drain_PE_8_9_V_full_n_pass_0_out),
    .fifo_cout_drain_PE_8_9_V_full_n_pass_1(fifo_cout_drain_PE_8_9_V_full_n_pass_1_in),
    .PE_wrapper255_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper255_U0_fifo_cout_drain_out_V_write_pass_0_in),
    .PE_wrapper255_U0_fifo_cout_drain_out_V_write_pass_1(PE_wrapper255_U0_fifo_cout_drain_out_V_write_pass_1_out),
    .PE_wrapper244_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper244_U0_fifo_w_out_V_V_din_pass_0_in),
    .PE_wrapper244_U0_fifo_w_out_V_V_din_pass_1(PE_wrapper244_U0_fifo_w_out_V_V_din_pass_1_out),
    .fifo_w_PE_7_11_V_V_full_n_pass_0(fifo_w_PE_7_11_V_V_full_n_pass_0_out),
    .fifo_w_PE_7_11_V_V_full_n_pass_1(fifo_w_PE_7_11_V_V_full_n_pass_1_in),
    .PE_wrapper244_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper244_U0_fifo_w_out_V_V_write_pass_0_in),
    .PE_wrapper244_U0_fifo_w_out_V_V_write_pass_1(PE_wrapper244_U0_fifo_w_out_V_V_write_pass_1_out),
    .cout_drain_IO_L1_out_wrapper517_U0_fifo_cout_drain_out_V_V_din_pass_1(cout_drain_IO_L1_out_wrapper517_U0_fifo_cout_drain_out_V_V_din_pass_1_in),
    .cout_drain_IO_L1_out_wrapper517_U0_fifo_cout_drain_out_V_V_din_pass_2(cout_drain_IO_L1_out_wrapper517_U0_fifo_cout_drain_out_V_V_din_pass_2_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_9_9_V_V_full_n_pass_1(fifo_cout_drain_cout_drain_IO_L1_out_9_9_V_V_full_n_pass_1_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_9_9_V_V_full_n_pass_2(fifo_cout_drain_cout_drain_IO_L1_out_9_9_V_V_full_n_pass_2_in),
    .cout_drain_IO_L1_out_wrapper517_U0_fifo_cout_drain_out_V_V_write_pass_1(cout_drain_IO_L1_out_wrapper517_U0_fifo_cout_drain_out_V_V_write_pass_1_in),
    .cout_drain_IO_L1_out_wrapper517_U0_fifo_cout_drain_out_V_V_write_pass_2(cout_drain_IO_L1_out_wrapper517_U0_fifo_cout_drain_out_V_V_write_pass_2_out),
    .PE_wrapper255_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper255_U0_fifo_w_out_V_V_din_pass_0_in),
    .PE_wrapper255_U0_fifo_w_out_V_V_din_pass_1(PE_wrapper255_U0_fifo_w_out_V_V_din_pass_1_out),
    .fifo_w_PE_8_10_V_V_full_n_pass_0(fifo_w_PE_8_10_V_V_full_n_pass_0_out),
    .fifo_w_PE_8_10_V_V_full_n_pass_1(fifo_w_PE_8_10_V_V_full_n_pass_1_in),
    .PE_wrapper255_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper255_U0_fifo_w_out_V_V_write_pass_0_in),
    .PE_wrapper255_U0_fifo_w_out_V_V_write_pass_1(PE_wrapper255_U0_fifo_w_out_V_V_write_pass_1_out),
    .PE_wrapper173_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper173_U0_fifo_cin_out_V_V_din_pass_0_in),
    .PE_wrapper173_U0_fifo_cin_out_V_V_din_pass_1(PE_wrapper173_U0_fifo_cin_out_V_V_din_pass_1_out),
    .fifo_cin_PE_2_11_V_V_full_n_pass_0(fifo_cin_PE_2_11_V_V_full_n_pass_0_out),
    .fifo_cin_PE_2_11_V_V_full_n_pass_1(fifo_cin_PE_2_11_V_V_full_n_pass_1_in),
    .PE_wrapper173_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper173_U0_fifo_cin_out_V_V_write_pass_0_in),
    .PE_wrapper173_U0_fifo_cin_out_V_V_write_pass_1(PE_wrapper173_U0_fifo_cin_out_V_V_write_pass_1_out),
    .cout_drain_IO_L1_out_wrapper533_U0_fifo_cout_drain_out_V_V_din_pass_1(cout_drain_IO_L1_out_wrapper533_U0_fifo_cout_drain_out_V_V_din_pass_1_in),
    .cout_drain_IO_L1_out_wrapper533_U0_fifo_cout_drain_out_V_V_din_pass_2(cout_drain_IO_L1_out_wrapper533_U0_fifo_cout_drain_out_V_V_din_pass_2_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_10_9_V_V_full_n_pass_1(fifo_cout_drain_cout_drain_IO_L1_out_10_9_V_V_full_n_pass_1_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_10_9_V_V_full_n_pass_2(fifo_cout_drain_cout_drain_IO_L1_out_10_9_V_V_full_n_pass_2_in),
    .cout_drain_IO_L1_out_wrapper533_U0_fifo_cout_drain_out_V_V_write_pass_1(cout_drain_IO_L1_out_wrapper533_U0_fifo_cout_drain_out_V_V_write_pass_1_in),
    .cout_drain_IO_L1_out_wrapper533_U0_fifo_cout_drain_out_V_V_write_pass_2(cout_drain_IO_L1_out_wrapper533_U0_fifo_cout_drain_out_V_V_write_pass_2_out),
    .PE_wrapper158_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper158_U0_fifo_w_out_V_V_din_pass_0_in),
    .fifo_w_PE_0_9_V_V_full_n_pass_0(fifo_w_PE_0_9_V_V_full_n_pass_0_out),
    .PE_wrapper158_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper158_U0_fifo_w_out_V_V_write_pass_0_in),
    .cout_drain_IO_L1_out_wrapper523_U0_fifo_cout_drain_out_V_V_din_pass_1(cout_drain_IO_L1_out_wrapper523_U0_fifo_cout_drain_out_V_V_din_pass_1_in),
    .fifo_cout_drain_cout_drain_IO_L1_out_9_3_V_V_full_n_pass_1(fifo_cout_drain_cout_drain_IO_L1_out_9_3_V_V_full_n_pass_1_out),
    .cout_drain_IO_L1_out_wrapper523_U0_fifo_cout_drain_out_V_V_write_pass_1(cout_drain_IO_L1_out_wrapper523_U0_fifo_cout_drain_out_V_V_write_pass_1_in),
    .PE_wrapper219_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper219_U0_fifo_w_out_V_V_din_pass_0_out),
    .fifo_w_PE_5_10_V_V_full_n_pass_0(fifo_w_PE_5_10_V_V_full_n_pass_0_in),
    .PE_wrapper219_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper219_U0_fifo_w_out_V_V_write_pass_0_out),
    .PE_wrapper170_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper170_U0_fifo_w_out_V_V_din_pass_0_in),
    .fifo_w_PE_1_9_V_V_full_n_pass_0(fifo_w_PE_1_9_V_V_full_n_pass_0_out),
    .PE_wrapper170_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper170_U0_fifo_w_out_V_V_write_pass_0_in),
    .PE_wrapper171_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper171_U0_fifo_cin_out_V_V_din_pass_0_out),
    .fifo_cin_PE_2_9_V_V_full_n_pass_0(fifo_cin_PE_2_9_V_V_full_n_pass_0_in),
    .PE_wrapper171_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper171_U0_fifo_cin_out_V_V_write_pass_0_out),
    .PE_wrapper172_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper172_U0_fifo_w_out_V_V_din_pass_0_out),
    .fifo_w_PE_1_11_V_V_full_n_pass_0(fifo_w_PE_1_11_V_V_full_n_pass_0_in),
    .PE_wrapper172_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper172_U0_fifo_w_out_V_V_write_pass_0_out),
    .cout_drain_IO_L2_out559_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L2_out559_U0_fifo_cout_drain_out_V_V_din_pass_0_out),
    .fifo_cout_drain_cout_drain_IO_L2_out_9_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L2_out_9_V_V_full_n_pass_0_in),
    .cout_drain_IO_L2_out559_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L2_out559_U0_fifo_cout_drain_out_V_V_write_pass_0_out),
    .PE_wrapper206_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper206_U0_fifo_w_out_V_V_din_pass_0_in),
    .fifo_w_PE_4_9_V_V_full_n_pass_0(fifo_w_PE_4_9_V_V_full_n_pass_0_out),
    .PE_wrapper206_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper206_U0_fifo_w_out_V_V_write_pass_0_in),
    .cin_IO_L2_in132_U0_fifo_cin_out_V_V_din_pass_0(cin_IO_L2_in132_U0_fifo_cin_out_V_V_din_pass_0_in),
    .fifo_cin_cin_IO_L2_in_9_V_V_full_n_pass_0(fifo_cin_cin_IO_L2_in_9_V_V_full_n_pass_0_out),
    .cin_IO_L2_in132_U0_fifo_cin_out_V_V_write_pass_0(cin_IO_L2_in132_U0_fifo_cin_out_V_V_write_pass_0_in),
    .PE_wrapper160_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper160_U0_fifo_w_out_V_V_din_pass_0_out),
    .fifo_w_PE_0_11_V_V_full_n_pass_0(fifo_w_PE_0_11_V_V_full_n_pass_0_in),
    .PE_wrapper160_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper160_U0_fifo_w_out_V_V_write_pass_0_out),
    .cout_drain_IO_L2_out558_U0_fifo_cout_drain_out_V_V_din_pass_1(cout_drain_IO_L2_out558_U0_fifo_cout_drain_out_V_V_din_pass_1_in),
    .fifo_cout_drain_cout_drain_IO_L2_out_10_V_V_full_n_pass_1(fifo_cout_drain_cout_drain_IO_L2_out_10_V_V_full_n_pass_1_out),
    .cout_drain_IO_L2_out558_U0_fifo_cout_drain_out_V_V_write_pass_1(cout_drain_IO_L2_out558_U0_fifo_cout_drain_out_V_V_write_pass_1_in),
    .PE_wrapper207_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper207_U0_fifo_w_out_V_V_din_pass_0_out),
    .fifo_w_PE_4_10_V_V_full_n_pass_0(fifo_w_PE_4_10_V_V_full_n_pass_0_in),
    .PE_wrapper207_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper207_U0_fifo_w_out_V_V_write_pass_0_out),
    .PE_wrapper183_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper183_U0_fifo_cout_drain_out_V_din_pass_0_in),
    .fifo_cout_drain_PE_2_9_V_full_n_pass_0(fifo_cout_drain_PE_2_9_V_full_n_pass_0_out),
    .PE_wrapper183_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper183_U0_fifo_cout_drain_out_V_write_pass_0_in),
    .cout_drain_IO_L1_out_wrapper522_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper522_U0_fifo_cout_drain_out_V_V_din_pass_0_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_9_4_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_9_4_V_V_full_n_pass_0_in),
    .cout_drain_IO_L1_out_wrapper522_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper522_U0_fifo_cout_drain_out_V_V_write_pass_0_out),
    .cout_drain_IO_L1_out_wrapper540_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper540_U0_fifo_cout_drain_out_V_V_din_pass_0_in),
    .fifo_cout_drain_cout_drain_IO_L1_out_10_2_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_10_2_V_V_full_n_pass_0_out),
    .cout_drain_IO_L1_out_wrapper540_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper540_U0_fifo_cout_drain_out_V_V_write_pass_0_in),
    .cout_drain_IO_L1_out_wrapper542_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper542_U0_fifo_cout_drain_out_V_V_din_pass_0_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_10_0_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_10_0_V_V_full_n_pass_0_in),
    .cout_drain_IO_L1_out_wrapper542_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper542_U0_fifo_cout_drain_out_V_V_write_pass_0_out),
    .PE_wrapper219_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper219_U0_fifo_cin_out_V_V_din_pass_0_out),
    .fifo_cin_PE_6_9_V_V_full_n_pass_0(fifo_cin_PE_6_9_V_V_full_n_pass_0_in),
    .PE_wrapper219_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper219_U0_fifo_cin_out_V_V_write_pass_0_out),
    .PE_wrapper172_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper172_U0_fifo_cin_out_V_V_din_pass_0_out),
    .fifo_cin_PE_2_10_V_V_full_n_pass_0(fifo_cin_PE_2_10_V_V_full_n_pass_0_in),
    .PE_wrapper172_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper172_U0_fifo_cin_out_V_V_write_pass_0_out),
    .PE_wrapper195_U0_fifo_cin_out_V_V_din_pass_1(PE_wrapper195_U0_fifo_cin_out_V_V_din_pass_1_in),
    .fifo_cin_PE_4_9_V_V_full_n_pass_1(fifo_cin_PE_4_9_V_V_full_n_pass_1_out),
    .PE_wrapper195_U0_fifo_cin_out_V_V_write_pass_1(PE_wrapper195_U0_fifo_cin_out_V_V_write_pass_1_in),
    .cin_IO_L2_in134_U0_fifo_cin_out_V_V_din_pass_0(cin_IO_L2_in134_U0_fifo_cin_out_V_V_din_pass_0_out),
    .fifo_cin_cin_IO_L2_in_11_V_V_full_n_pass_0(fifo_cin_cin_IO_L2_in_11_V_V_full_n_pass_0_in),
    .cin_IO_L2_in134_U0_fifo_cin_out_V_V_write_pass_0(cin_IO_L2_in134_U0_fifo_cin_out_V_V_write_pass_0_out),
    .PE_wrapper218_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper218_U0_fifo_w_out_V_V_din_pass_0_in),
    .fifo_w_PE_5_9_V_V_full_n_pass_0(fifo_w_PE_5_9_V_V_full_n_pass_0_out),
    .PE_wrapper218_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper218_U0_fifo_w_out_V_V_write_pass_0_in),
    .cout_drain_IO_L1_out_wrapper521_U0_fifo_cout_drain_out_V_V_din_pass_1(cout_drain_IO_L1_out_wrapper521_U0_fifo_cout_drain_out_V_V_din_pass_1_in),
    .fifo_cout_drain_cout_drain_IO_L1_out_9_5_V_V_full_n_pass_1(fifo_cout_drain_cout_drain_IO_L1_out_9_5_V_V_full_n_pass_1_out),
    .cout_drain_IO_L1_out_wrapper521_U0_fifo_cout_drain_out_V_V_write_pass_1(cout_drain_IO_L1_out_wrapper521_U0_fifo_cout_drain_out_V_V_write_pass_1_in),
    .PE_wrapper219_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper219_U0_fifo_cout_drain_out_V_din_pass_0_out),
    .fifo_cout_drain_PE_5_9_V_full_n_pass_0(fifo_cout_drain_PE_5_9_V_full_n_pass_0_in),
    .PE_wrapper219_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper219_U0_fifo_cout_drain_out_V_write_pass_0_out),
    .ap_clk(ap_clk),
    .ap_start_Boundary_X6Y12_To_X8Y12(ap_start_Boundary_X6Y12_To_X8Y12_in),
    .ap_rst_n_Boundary_X6Y12_To_X8Y12(ap_rst_n_Boundary_X6Y12_To_X8Y12_in),
    .ap_done_Boundary_X6Y12_To_X8Y12(ap_done_Boundary_X6Y12_To_X8Y12_out),
    .ap_start_Boundary_X6Y14_To_X8Y14(ap_start_Boundary_X6Y14_To_X8Y14_out),
    .ap_rst_n_Boundary_X6Y14_To_X8Y14(ap_rst_n_Boundary_X6Y14_To_X8Y14_out),
    .ap_done_Boundary_X6Y14_To_X8Y14(ap_done_Boundary_X6Y14_To_X8Y14_in)
  );


  (* keep_hierarchy = "yes" *) CR_X6Y14_To_CR_X7Y15_ctrl CR_X6Y14_To_CR_X7Y15_ctrl_U0 (
    .PE_wrapper231_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper231_U0_fifo_cin_out_V_V_din_pass_0_in),
    .PE_wrapper231_U0_fifo_cin_out_V_V_din_pass_1(PE_wrapper231_U0_fifo_cin_out_V_V_din_pass_1_out),
    .fifo_cin_PE_7_9_V_V_full_n_pass_0(fifo_cin_PE_7_9_V_V_full_n_pass_0_out),
    .fifo_cin_PE_7_9_V_V_full_n_pass_1(fifo_cin_PE_7_9_V_V_full_n_pass_1_in),
    .PE_wrapper231_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper231_U0_fifo_cin_out_V_V_write_pass_0_in),
    .PE_wrapper231_U0_fifo_cin_out_V_V_write_pass_1(PE_wrapper231_U0_fifo_cin_out_V_V_write_pass_1_out),
    .cout_drain_IO_L1_out_wrapper523_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper523_U0_fifo_cout_drain_out_V_V_din_pass_0_in),
    .cout_drain_IO_L1_out_wrapper523_U0_fifo_cout_drain_out_V_V_din_pass_1(cout_drain_IO_L1_out_wrapper523_U0_fifo_cout_drain_out_V_V_din_pass_1_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_9_3_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_9_3_V_V_full_n_pass_0_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_9_3_V_V_full_n_pass_1(fifo_cout_drain_cout_drain_IO_L1_out_9_3_V_V_full_n_pass_1_in),
    .cout_drain_IO_L1_out_wrapper523_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper523_U0_fifo_cout_drain_out_V_V_write_pass_0_in),
    .cout_drain_IO_L1_out_wrapper523_U0_fifo_cout_drain_out_V_V_write_pass_1(cout_drain_IO_L1_out_wrapper523_U0_fifo_cout_drain_out_V_V_write_pass_1_out),
    .cout_drain_IO_L2_out558_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L2_out558_U0_fifo_cout_drain_out_V_V_din_pass_0_in),
    .cout_drain_IO_L2_out558_U0_fifo_cout_drain_out_V_V_din_pass_1(cout_drain_IO_L2_out558_U0_fifo_cout_drain_out_V_V_din_pass_1_out),
    .fifo_cout_drain_cout_drain_IO_L2_out_10_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L2_out_10_V_V_full_n_pass_0_out),
    .fifo_cout_drain_cout_drain_IO_L2_out_10_V_V_full_n_pass_1(fifo_cout_drain_cout_drain_IO_L2_out_10_V_V_full_n_pass_1_in),
    .cout_drain_IO_L2_out558_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L2_out558_U0_fifo_cout_drain_out_V_V_write_pass_0_in),
    .cout_drain_IO_L2_out558_U0_fifo_cout_drain_out_V_V_write_pass_1(cout_drain_IO_L2_out558_U0_fifo_cout_drain_out_V_V_write_pass_1_out),
    .PE_wrapper195_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper195_U0_fifo_cin_out_V_V_din_pass_0_in),
    .PE_wrapper195_U0_fifo_cin_out_V_V_din_pass_1(PE_wrapper195_U0_fifo_cin_out_V_V_din_pass_1_out),
    .fifo_cin_PE_4_9_V_V_full_n_pass_0(fifo_cin_PE_4_9_V_V_full_n_pass_0_out),
    .fifo_cin_PE_4_9_V_V_full_n_pass_1(fifo_cin_PE_4_9_V_V_full_n_pass_1_in),
    .PE_wrapper195_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper195_U0_fifo_cin_out_V_V_write_pass_0_in),
    .PE_wrapper195_U0_fifo_cin_out_V_V_write_pass_1(PE_wrapper195_U0_fifo_cin_out_V_V_write_pass_1_out),
    .cout_drain_IO_L1_out_wrapper521_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper521_U0_fifo_cout_drain_out_V_V_din_pass_0_in),
    .cout_drain_IO_L1_out_wrapper521_U0_fifo_cout_drain_out_V_V_din_pass_1(cout_drain_IO_L1_out_wrapper521_U0_fifo_cout_drain_out_V_V_din_pass_1_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_9_5_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_9_5_V_V_full_n_pass_0_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_9_5_V_V_full_n_pass_1(fifo_cout_drain_cout_drain_IO_L1_out_9_5_V_V_full_n_pass_1_in),
    .cout_drain_IO_L1_out_wrapper521_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper521_U0_fifo_cout_drain_out_V_V_write_pass_0_in),
    .cout_drain_IO_L1_out_wrapper521_U0_fifo_cout_drain_out_V_V_write_pass_1(cout_drain_IO_L1_out_wrapper521_U0_fifo_cout_drain_out_V_V_write_pass_1_out),
    .cout_drain_IO_L1_out_wrapper551_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper551_U0_fifo_cout_drain_out_V_V_din_pass_0_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_11_6_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_11_6_V_V_full_n_pass_0_in),
    .cout_drain_IO_L1_out_wrapper551_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper551_U0_fifo_cout_drain_out_V_V_write_pass_0_out),
    .cout_drain_IO_L1_out_wrapper556_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper556_U0_fifo_cout_drain_out_V_V_din_pass_0_in),
    .fifo_cout_drain_cout_drain_IO_L1_out_11_1_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_11_1_V_V_full_n_pass_0_out),
    .cout_drain_IO_L1_out_wrapper556_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper556_U0_fifo_cout_drain_out_V_V_write_pass_0_in),
    .PE_wrapper160_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper160_U0_fifo_w_out_V_V_din_pass_0_in),
    .fifo_w_PE_0_11_V_V_full_n_pass_0(fifo_w_PE_0_11_V_V_full_n_pass_0_out),
    .PE_wrapper160_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper160_U0_fifo_w_out_V_V_write_pass_0_in),
    .PE_wrapper244_U0_fifo_cin_out_V_V_din_pass_1(PE_wrapper244_U0_fifo_cin_out_V_V_din_pass_1_in),
    .fifo_cin_PE_8_10_V_V_full_n_pass_1(fifo_cin_PE_8_10_V_V_full_n_pass_1_out),
    .PE_wrapper244_U0_fifo_cin_out_V_V_write_pass_1(PE_wrapper244_U0_fifo_cin_out_V_V_write_pass_1_in),
    .PE_wrapper173_U0_fifo_w_out_V_V_din_pass_1(PE_wrapper173_U0_fifo_w_out_V_V_din_pass_1_in),
    .fifo_w_PE_1_12_V_V_full_n_pass_1(fifo_w_PE_1_12_V_V_full_n_pass_1_out),
    .PE_wrapper173_U0_fifo_w_out_V_V_write_pass_1(PE_wrapper173_U0_fifo_w_out_V_V_write_pass_1_in),
    .PE_wrapper184_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper184_U0_fifo_w_out_V_V_din_pass_0_in),
    .fifo_w_PE_2_11_V_V_full_n_pass_0(fifo_w_PE_2_11_V_V_full_n_pass_0_out),
    .PE_wrapper184_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper184_U0_fifo_w_out_V_V_write_pass_0_in),
    .PE_wrapper161_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper161_U0_fifo_cin_out_V_V_din_pass_0_out),
    .fifo_cin_PE_1_11_V_V_full_n_pass_0(fifo_cin_PE_1_11_V_V_full_n_pass_0_in),
    .PE_wrapper161_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper161_U0_fifo_cin_out_V_V_write_pass_0_out),
    .PE_wrapper256_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper256_U0_fifo_cin_out_V_V_din_pass_0_out),
    .fifo_cin_PE_9_10_V_V_full_n_pass_0(fifo_cin_PE_9_10_V_V_full_n_pass_0_in),
    .PE_wrapper256_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper256_U0_fifo_cin_out_V_V_write_pass_0_out),
    .PE_wrapper196_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper196_U0_fifo_w_out_V_V_din_pass_0_in),
    .fifo_w_PE_3_11_V_V_full_n_pass_0(fifo_w_PE_3_11_V_V_full_n_pass_0_out),
    .PE_wrapper196_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper196_U0_fifo_w_out_V_V_write_pass_0_in),
    .PE_wrapper209_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper209_U0_fifo_w_out_V_V_din_pass_0_in),
    .fifo_w_PE_4_12_V_V_full_n_pass_0(fifo_w_PE_4_12_V_V_full_n_pass_0_out),
    .PE_wrapper209_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper209_U0_fifo_w_out_V_V_write_pass_0_in),
    .PE_wrapper233_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper233_U0_fifo_cin_out_V_V_din_pass_0_in),
    .fifo_cin_PE_7_11_V_V_full_n_pass_0(fifo_cin_PE_7_11_V_V_full_n_pass_0_out),
    .PE_wrapper233_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper233_U0_fifo_cin_out_V_V_write_pass_0_in),
    .PE_wrapper255_U0_fifo_cout_drain_out_V_din_pass_1(PE_wrapper255_U0_fifo_cout_drain_out_V_din_pass_1_in),
    .fifo_cout_drain_PE_8_9_V_full_n_pass_1(fifo_cout_drain_PE_8_9_V_full_n_pass_1_out),
    .PE_wrapper255_U0_fifo_cout_drain_out_V_write_pass_1(PE_wrapper255_U0_fifo_cout_drain_out_V_write_pass_1_in),
    .PE_wrapper197_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper197_U0_fifo_cin_out_V_V_din_pass_0_out),
    .fifo_cin_PE_4_11_V_V_full_n_pass_0(fifo_cin_PE_4_11_V_V_full_n_pass_0_in),
    .PE_wrapper197_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper197_U0_fifo_cin_out_V_V_write_pass_0_out),
    .PE_wrapper185_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper185_U0_fifo_cout_drain_out_V_din_pass_0_out),
    .fifo_cout_drain_PE_2_11_V_full_n_pass_0(fifo_cout_drain_PE_2_11_V_full_n_pass_0_in),
    .PE_wrapper185_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper185_U0_fifo_cout_drain_out_V_write_pass_0_out),
    .cout_drain_IO_L1_out_wrapper518_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper518_U0_fifo_cout_drain_out_V_V_din_pass_0_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_9_8_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_9_8_V_V_full_n_pass_0_in),
    .cout_drain_IO_L1_out_wrapper518_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper518_U0_fifo_cout_drain_out_V_V_write_pass_0_out),
    .PE_wrapper244_U0_fifo_w_out_V_V_din_pass_1(PE_wrapper244_U0_fifo_w_out_V_V_din_pass_1_in),
    .fifo_w_PE_7_11_V_V_full_n_pass_1(fifo_w_PE_7_11_V_V_full_n_pass_1_out),
    .PE_wrapper244_U0_fifo_w_out_V_V_write_pass_1(PE_wrapper244_U0_fifo_w_out_V_V_write_pass_1_in),
    .cout_drain_IO_L1_out_wrapper517_U0_fifo_cout_drain_out_V_V_din_pass_2(cout_drain_IO_L1_out_wrapper517_U0_fifo_cout_drain_out_V_V_din_pass_2_in),
    .fifo_cout_drain_cout_drain_IO_L1_out_9_9_V_V_full_n_pass_2(fifo_cout_drain_cout_drain_IO_L1_out_9_9_V_V_full_n_pass_2_out),
    .cout_drain_IO_L1_out_wrapper517_U0_fifo_cout_drain_out_V_V_write_pass_2(cout_drain_IO_L1_out_wrapper517_U0_fifo_cout_drain_out_V_V_write_pass_2_in),
    .cout_drain_IO_L1_out_wrapper549_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper549_U0_fifo_cout_drain_out_V_V_din_pass_0_in),
    .fifo_cout_drain_cout_drain_IO_L1_out_11_8_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_11_8_V_V_full_n_pass_0_out),
    .cout_drain_IO_L1_out_wrapper549_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper549_U0_fifo_cout_drain_out_V_V_write_pass_0_in),
    .PE_wrapper255_U0_fifo_w_out_V_V_din_pass_1(PE_wrapper255_U0_fifo_w_out_V_V_din_pass_1_in),
    .fifo_w_PE_8_10_V_V_full_n_pass_1(fifo_w_PE_8_10_V_V_full_n_pass_1_out),
    .PE_wrapper255_U0_fifo_w_out_V_V_write_pass_1(PE_wrapper255_U0_fifo_w_out_V_V_write_pass_1_in),
    .cout_drain_IO_L1_out_wrapper534_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper534_U0_fifo_cout_drain_out_V_V_din_pass_0_out),
    .fifo_cout_drain_cout_drain_IO_L1_out_10_8_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_10_8_V_V_full_n_pass_0_in),
    .cout_drain_IO_L1_out_wrapper534_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper534_U0_fifo_cout_drain_out_V_V_write_pass_0_out),
    .PE_wrapper257_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper257_U0_fifo_cin_out_V_V_din_pass_0_out),
    .fifo_cin_PE_9_11_V_V_full_n_pass_0(fifo_cin_PE_9_11_V_V_full_n_pass_0_in),
    .PE_wrapper257_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper257_U0_fifo_cin_out_V_V_write_pass_0_out),
    .PE_wrapper257_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper257_U0_fifo_cout_drain_out_V_din_pass_0_out),
    .fifo_cout_drain_PE_8_11_V_full_n_pass_0(fifo_cout_drain_PE_8_11_V_full_n_pass_0_in),
    .PE_wrapper257_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper257_U0_fifo_cout_drain_out_V_write_pass_0_out),
    .cin_IO_L2_in_boundary_U0_fifo_cin_local_out_V_V_din_pass_0(cin_IO_L2_in_boundary_U0_fifo_cin_local_out_V_V_din_pass_0_in),
    .fifo_cin_PE_0_11_V_V_full_n_pass_0(fifo_cin_PE_0_11_V_V_full_n_pass_0_out),
    .cin_IO_L2_in_boundary_U0_fifo_cin_local_out_V_V_write_pass_0(cin_IO_L2_in_boundary_U0_fifo_cin_local_out_V_V_write_pass_0_in),
    .PE_wrapper173_U0_fifo_cin_out_V_V_din_pass_1(PE_wrapper173_U0_fifo_cin_out_V_V_din_pass_1_in),
    .fifo_cin_PE_2_11_V_V_full_n_pass_1(fifo_cin_PE_2_11_V_V_full_n_pass_1_out),
    .PE_wrapper173_U0_fifo_cin_out_V_V_write_pass_1(PE_wrapper173_U0_fifo_cin_out_V_V_write_pass_1_in),
    .cout_drain_IO_L1_out_wrapper533_U0_fifo_cout_drain_out_V_V_din_pass_2(cout_drain_IO_L1_out_wrapper533_U0_fifo_cout_drain_out_V_V_din_pass_2_in),
    .fifo_cout_drain_cout_drain_IO_L1_out_10_9_V_V_full_n_pass_2(fifo_cout_drain_cout_drain_IO_L1_out_10_9_V_V_full_n_pass_2_out),
    .cout_drain_IO_L1_out_wrapper533_U0_fifo_cout_drain_out_V_V_write_pass_2(cout_drain_IO_L1_out_wrapper533_U0_fifo_cout_drain_out_V_V_write_pass_2_in),
    .PE_wrapper197_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper197_U0_fifo_cout_drain_out_V_din_pass_0_out),
    .fifo_cout_drain_PE_3_11_V_full_n_pass_0(fifo_cout_drain_PE_3_11_V_full_n_pass_0_in),
    .PE_wrapper197_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper197_U0_fifo_cout_drain_out_V_write_pass_0_out),
    .PE_wrapper233_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper233_U0_fifo_cout_drain_out_V_din_pass_0_in),
    .fifo_cout_drain_PE_6_11_V_full_n_pass_0(fifo_cout_drain_PE_6_11_V_full_n_pass_0_out),
    .PE_wrapper233_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper233_U0_fifo_cout_drain_out_V_write_pass_0_in),
    .PE_wrapper185_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper185_U0_fifo_w_out_V_V_din_pass_0_out),
    .fifo_w_PE_2_12_V_V_full_n_pass_0(fifo_w_PE_2_12_V_V_full_n_pass_0_in),
    .PE_wrapper185_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper185_U0_fifo_w_out_V_V_write_pass_0_out),
    .cout_drain_IO_L2_out_boundary_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L2_out_boundary_U0_fifo_cout_drain_out_V_V_din_pass_0_out),
    .fifo_cout_drain_cout_drain_IO_L2_out_11_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L2_out_11_V_V_full_n_pass_0_in),
    .cout_drain_IO_L2_out_boundary_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L2_out_boundary_U0_fifo_cout_drain_out_V_V_write_pass_0_out),
    .ap_clk(ap_clk),
    .ap_start_Boundary_X6Y14_To_X8Y14(ap_start_Boundary_X6Y14_To_X8Y14_in),
    .ap_rst_n_Boundary_X6Y14_To_X8Y14(ap_rst_n_Boundary_X6Y14_To_X8Y14_in),
    .ap_done_Boundary_X6Y14_To_X8Y14(ap_done_Boundary_X6Y14_To_X8Y14_out)
  );
endmodule

// first-word fall-through (FWFT) FIFO
// if its capacity > THRESHOLD bits, it uses block RAM, otherwise it will uses
// shift register LUT
module fifo_almost_full #(
  parameter DATA_WIDTH = 32,
  parameter ADDR_WIDTH = 5,
  parameter DEPTH      = 32,
  parameter THRESHOLD  = 18432,
  parameter GRACE_PERIOD = 2
) (
  input wire clk,
  input wire reset,
  // write
  output wire                  if_full_n,
  input  wire                  if_write_ce,
  input  wire                  if_write,
  input  wire [DATA_WIDTH-1:0] if_din,
  // read
  output wire                  if_empty_n,
  input  wire                  if_read_ce,
  input  wire                  if_read,
  output wire [DATA_WIDTH-1:0] if_dout
);
  parameter REAL_DEPTH = GRACE_PERIOD + DEPTH + 4;
  parameter REAL_ADDR_WIDTH  = $clog2(REAL_DEPTH);
generate
  if (DATA_WIDTH * DEPTH > THRESHOLD) begin : bram
    fifo_bram_almost_full #(
      .DATA_WIDTH(DATA_WIDTH),
      .ADDR_WIDTH(REAL_ADDR_WIDTH),
      .DEPTH     (REAL_DEPTH),
      .GRACE_PERIOD(GRACE_PERIOD) /*********/
    ) unit (
      .clk  (clk),
      .reset(reset),
      .if_full_n  (if_full_n),
      .if_write_ce(if_write_ce),
      .if_write   (if_write),
      .if_din     (if_din),
      .if_empty_n(if_empty_n),
      .if_read_ce(if_read_ce),
      .if_read   (if_read),
      .if_dout   (if_dout)
    );
  end else begin : srl
    fifo_srl_almost_full #(
      .DATA_WIDTH(DATA_WIDTH),
      .ADDR_WIDTH(REAL_ADDR_WIDTH),
      .DEPTH     (REAL_DEPTH),
      .GRACE_PERIOD(GRACE_PERIOD) /*********/
    ) unit (
      .clk  (clk),
      .reset(reset),
      .if_full_n  (if_full_n),
      .if_write_ce(if_write_ce),
      .if_write   (if_write),
      .if_din     (if_din),
      .if_empty_n(if_empty_n),
      .if_read_ce(if_read_ce),
      .if_read   (if_read),
      .if_dout   (if_dout)
    );
  end
endgenerate
endmodule  // fifo
/////////////////////////////////////////////////////////////////
module fifo_srl_almost_full (
    clk,
    reset,
    if_empty_n,
    if_read_ce,
    if_read,
    if_dout,
    if_full_n,
    if_write_ce,
    if_write,
    if_din);
parameter MEM_STYLE   = "shiftreg";
parameter DATA_WIDTH  = 32'd32;
parameter ADDR_WIDTH  = 32'd4;
parameter DEPTH       = 5'd16;
/*******************************************/
parameter GRACE_PERIOD = 2;
/*******************************************/
input clk;
input reset;
output if_empty_n;
input if_read_ce;
input if_read;
output[DATA_WIDTH - 1:0] if_dout;
output if_full_n;
input if_write_ce;
input if_write;
input[DATA_WIDTH - 1:0] if_din;
wire[ADDR_WIDTH - 1:0] shiftReg_addr ;
wire[DATA_WIDTH - 1:0] shiftReg_data, shiftReg_q;
wire                     shiftReg_ce;
reg[ADDR_WIDTH:0] mOutPtr = ~{(ADDR_WIDTH+1){1'b0}};
reg internal_empty_n = 0, internal_full_n = 1;
assign if_empty_n = internal_empty_n;
/*******************************************/
// assign if_full_n = internal_full_n;
wire almost_full = mOutPtr >= DEPTH - 1 - GRACE_PERIOD && mOutPtr != ~{ADDR_WIDTH+1{1'b0}};
assign if_full_n = ~almost_full;
/*******************************************/
assign shiftReg_data = if_din;
assign if_dout = shiftReg_q;
always @ (posedge clk) begin
    if (reset == 1'b1)
    begin
        mOutPtr <= ~{ADDR_WIDTH+1{1'b0}};
        internal_empty_n <= 1'b0;
        internal_full_n <= 1'b1;
    end
    else begin
        if (((if_read & if_read_ce) == 1 & internal_empty_n == 1) && 
            ((if_write & if_write_ce) == 0 | internal_full_n == 0))
        begin
            mOutPtr <= mOutPtr - 5'd1;
            if (mOutPtr == 0)
                internal_empty_n <= 1'b0;
            internal_full_n <= 1'b1;
        end 
        else if (((if_read & if_read_ce) == 0 | internal_empty_n == 0) && 
            ((if_write & if_write_ce) == 1 & internal_full_n == 1))
        begin
            mOutPtr <= mOutPtr + 5'd1;
            internal_empty_n <= 1'b1;
            if (mOutPtr == DEPTH - 5'd2)
                internal_full_n <= 1'b0;
        end 
    end
end
assign shiftReg_addr = mOutPtr[ADDR_WIDTH] == 1'b0 ? mOutPtr[ADDR_WIDTH-1:0]:{ADDR_WIDTH{1'b0}};
assign shiftReg_ce = (if_write & if_write_ce) & internal_full_n;
fifo_srl_almost_full_internal 
#(
    .DATA_WIDTH(DATA_WIDTH),
    .ADDR_WIDTH(ADDR_WIDTH),
    .DEPTH(DEPTH))
U_fifo_w32_d16_A_ram (
    .clk(clk),
    .data(shiftReg_data),
    .ce(shiftReg_ce),
    .a(shiftReg_addr),
    .q(shiftReg_q));
endmodule  
module fifo_srl_almost_full_internal (
    clk,
    data,
    ce,
    a,
    q);
parameter DATA_WIDTH = 32'd32;
parameter ADDR_WIDTH = 32'd4;
parameter DEPTH = 5'd16;
input clk;
input [DATA_WIDTH-1:0] data;
input ce;
input [ADDR_WIDTH-1:0] a;
output [DATA_WIDTH-1:0] q;
reg[DATA_WIDTH-1:0] SRL_SIG [0:DEPTH-1];
integer i;
always @ (posedge clk)
    begin
        if (ce)
        begin
            for (i=0;i<DEPTH-1;i=i+1)
                SRL_SIG[i+1] <= SRL_SIG[i];
            SRL_SIG[0] <= data;
        end
    end
assign q = SRL_SIG[a];
endmodule
///////////////////////////////////////////////////////////
// first-word fall-through (FWFT) FIFO using block RAM or URAM (let Vivado choose)
// based on HLS generated code
module fifo_bram_almost_full #(
  parameter MEM_STYLE  = "auto",
  parameter DATA_WIDTH = 32,
  parameter ADDR_WIDTH = 5,
  parameter DEPTH      = 32,
  parameter GRACE_PERIOD = 2
) (
  input wire clk,
  input wire reset,
  // write
  output wire                  if_full_n,
  input  wire                  if_write_ce,
  input  wire                  if_write,
  input  wire [DATA_WIDTH-1:0] if_din,
  // read
  output wire                  if_empty_n,
  input  wire                  if_read_ce,
  input  wire                  if_read,
  output wire [DATA_WIDTH-1:0] if_dout
);
(* ram_style = MEM_STYLE *)
reg  [DATA_WIDTH-1:0] mem[0:DEPTH-1];
reg  [DATA_WIDTH-1:0] q_buf;
reg  [ADDR_WIDTH-1:0] waddr;
reg  [ADDR_WIDTH-1:0] raddr;
wire [ADDR_WIDTH-1:0] wnext;
wire [ADDR_WIDTH-1:0] rnext;
wire                  push;
wire                  pop;
reg  [ADDR_WIDTH-1:0] used;
reg                   full_n;
reg                   empty_n;
reg  [DATA_WIDTH-1:0] q_tmp;
reg                   show_ahead;
reg  [DATA_WIDTH-1:0] dout_buf;
reg                   dout_valid;
localparam DepthM1 = DEPTH[ADDR_WIDTH-1:0] - 1'd1;
/**************************************/
wire almost_full = (used >= DEPTH - 1 - GRACE_PERIOD);
//assign if_full_n  = full_n;
assign if_full_n  = ~almost_full;
/**************************************/
assign if_empty_n = dout_valid;
assign if_dout    = dout_buf;
assign push       = full_n & if_write_ce & if_write;
assign pop        = empty_n & if_read_ce & (~dout_valid | if_read);
assign wnext      = !push              ? waddr              :
                    (waddr == DepthM1) ? {ADDR_WIDTH{1'b0}} : waddr + 1'd1;
assign rnext      = !pop               ? raddr              :
                    (raddr == DepthM1) ? {ADDR_WIDTH{1'b0}} : raddr + 1'd1;
// waddr
always @(posedge clk) begin
  if (reset)
    waddr <= {ADDR_WIDTH{1'b0}};
  else
    waddr <= wnext;
end
// raddr
always @(posedge clk) begin
  if (reset)
    raddr <= {ADDR_WIDTH{1'b0}};
  else
    raddr <= rnext;
end
// used
always @(posedge clk) begin
  if (reset)
    used <= {ADDR_WIDTH{1'b0}};
  else if (push && !pop)
    used <= used + 1'b1;
  else if (!push && pop)
    used <= used - 1'b1;
end
// full_n
always @(posedge clk) begin
  if (reset)
    full_n <= 1'b1;
  else if (push && !pop)
    full_n <= (used != DepthM1);
  else if (!push && pop)
    full_n <= 1'b1;
end
// empty_n
always @(posedge clk) begin
  if (reset)
    empty_n <= 1'b0;
  else if (push && !pop)
    empty_n <= 1'b1;
  else if (!push && pop)
    empty_n <= (used != {{(ADDR_WIDTH-1){1'b0}},1'b1});
end
// mem
always @(posedge clk) begin
  if (push)
    mem[waddr] <= if_din;
end
// q_buf
always @(posedge clk) begin
  q_buf <= mem[rnext];
end
// q_tmp
always @(posedge clk) begin
  if (reset)
    q_tmp <= {DATA_WIDTH{1'b0}};
  else if (push)
    q_tmp <= if_din;
end
// show_ahead
always @(posedge clk) begin
  if (reset)
    show_ahead <= 1'b0;
  else if (push && used == {{(ADDR_WIDTH-1){1'b0}},pop})
    show_ahead <= 1'b1;
  else
    show_ahead <= 1'b0;
end
// dout_buf
always @(posedge clk) begin
  if (reset)
    dout_buf <= {DATA_WIDTH{1'b0}};
  else if (pop)
    dout_buf <= show_ahead? q_tmp : q_buf;
end
// dout_valid
always @(posedge clk) begin
  if (reset)
    dout_valid <= 1'b0;
  else if (pop)
    dout_valid <= 1'b1;
  else if (if_read_ce & if_read)
    dout_valid <= 1'b0;
end
endmodule  // fifo_bram

