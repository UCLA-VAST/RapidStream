

`timescale 1 ns / 1 ps
module CR_X4Y12_To_CR_X5Y13 (
  cout_drain_IO_L1_out_wrapper535_U0_fifo_cout_drain_out_V_V_din,
  fifo_cout_drain_cout_drain_IO_L1_out_10_7_V_V_full_n,
  cout_drain_IO_L1_out_wrapper535_U0_fifo_cout_drain_out_V_V_write,
  PE_wrapper219_U0_fifo_w_out_V_V_din,
  fifo_w_PE_5_10_V_V_full_n,
  PE_wrapper219_U0_fifo_w_out_V_V_write,
  cout_drain_IO_L1_out_wrapper537_U0_fifo_cout_drain_out_V_V_din,
  fifo_cout_drain_cout_drain_IO_L1_out_10_5_V_V_full_n,
  cout_drain_IO_L1_out_wrapper537_U0_fifo_cout_drain_out_V_V_write,
  PE_wrapper171_U0_fifo_cin_out_V_V_din,
  fifo_cin_PE_2_9_V_V_full_n,
  PE_wrapper171_U0_fifo_cin_out_V_V_write,
  PE_wrapper172_U0_fifo_w_out_V_V_din,
  fifo_w_PE_1_11_V_V_full_n,
  PE_wrapper172_U0_fifo_w_out_V_V_write,
  cout_drain_IO_L1_out_wrapper551_U0_fifo_cout_drain_out_V_V_din,
  fifo_cout_drain_cout_drain_IO_L1_out_11_6_V_V_full_n,
  cout_drain_IO_L1_out_wrapper551_U0_fifo_cout_drain_out_V_V_write,
  cout_drain_IO_L1_out_wrapper555_U0_fifo_cout_drain_out_V_V_din,
  fifo_cout_drain_cout_drain_IO_L1_out_11_2_V_V_full_n,
  cout_drain_IO_L1_out_wrapper555_U0_fifo_cout_drain_out_V_V_write,
  PE_wrapper196_U0_fifo_cin_out_V_V_din,
  fifo_cin_PE_4_10_V_V_full_n,
  PE_wrapper196_U0_fifo_cin_out_V_V_write,
  cout_drain_IO_L1_out_wrapper539_U0_fifo_cout_drain_out_V_V_din,
  fifo_cout_drain_cout_drain_IO_L1_out_10_3_V_V_full_n,
  cout_drain_IO_L1_out_wrapper539_U0_fifo_cout_drain_out_V_V_write,
  PE_wrapper244_U0_fifo_cin_out_V_V_din,
  fifo_cin_PE_8_10_V_V_full_n,
  PE_wrapper244_U0_fifo_cin_out_V_V_write,
  PE_wrapper231_U0_fifo_w_out_V_V_din,
  fifo_w_PE_6_10_V_V_full_n,
  PE_wrapper231_U0_fifo_w_out_V_V_write,
  PE_wrapper173_U0_fifo_w_out_V_V_din,
  fifo_w_PE_1_12_V_V_full_n,
  PE_wrapper173_U0_fifo_w_out_V_V_write,
  PE_wrapper231_U0_fifo_cout_drain_out_V_din,
  fifo_cout_drain_PE_6_9_V_full_n,
  PE_wrapper231_U0_fifo_cout_drain_out_V_write,
  PE_wrapper207_U0_fifo_w_out_V_V_din,
  fifo_w_PE_4_10_V_V_full_n,
  PE_wrapper207_U0_fifo_w_out_V_V_write,
  PE_wrapper221_U0_fifo_cout_drain_out_V_din,
  fifo_cout_drain_PE_5_11_V_full_n,
  PE_wrapper221_U0_fifo_cout_drain_out_V_write,
  PE_wrapper183_U0_fifo_cout_drain_out_V_din,
  fifo_cout_drain_PE_2_9_V_full_n,
  PE_wrapper183_U0_fifo_cout_drain_out_V_write,
  PE_wrapper161_U0_fifo_cin_out_V_V_din,
  fifo_cin_PE_1_11_V_V_full_n,
  PE_wrapper161_U0_fifo_cin_out_V_V_write,
  PE_wrapper232_U0_fifo_cout_drain_out_V_din,
  fifo_cout_drain_PE_6_10_V_full_n,
  PE_wrapper232_U0_fifo_cout_drain_out_V_write,
  kernel0_entry12_U0_cout_V_out_din,
  cout_V_c_full_n,
  kernel0_entry12_U0_cout_V_out_write,
  cout_drain_IO_L1_out_wrapper540_U0_fifo_cout_drain_out_V_V_din,
  fifo_cout_drain_cout_drain_IO_L1_out_10_2_V_V_full_n,
  cout_drain_IO_L1_out_wrapper540_U0_fifo_cout_drain_out_V_V_write,
  cout_drain_IO_L1_out_wrapper552_U0_fifo_cout_drain_out_V_V_din,
  fifo_cout_drain_cout_drain_IO_L1_out_11_5_V_V_full_n,
  cout_drain_IO_L1_out_wrapper552_U0_fifo_cout_drain_out_V_V_write,
  PE_wrapper243_U0_fifo_w_out_V_V_din,
  fifo_w_PE_7_10_V_V_full_n,
  PE_wrapper243_U0_fifo_w_out_V_V_write,
  PE_wrapper243_U0_fifo_cout_drain_out_V_din,
  fifo_cout_drain_PE_7_9_V_full_n,
  PE_wrapper243_U0_fifo_cout_drain_out_V_write,
  PE_wrapper184_U0_fifo_cout_drain_out_V_din,
  fifo_cout_drain_PE_2_10_V_full_n,
  PE_wrapper184_U0_fifo_cout_drain_out_V_write,
  PE_wrapper243_U0_fifo_cin_out_V_V_din,
  fifo_cin_PE_8_9_V_V_full_n,
  PE_wrapper243_U0_fifo_cin_out_V_V_write,
  PE_wrapper255_U0_fifo_cout_drain_out_V_din,
  fifo_cout_drain_PE_8_9_V_full_n,
  PE_wrapper255_U0_fifo_cout_drain_out_V_write,
  PE_wrapper185_U0_fifo_cout_drain_out_V_din,
  fifo_cout_drain_PE_2_11_V_full_n,
  PE_wrapper185_U0_fifo_cout_drain_out_V_write,
  cout_drain_IO_L1_out_wrapper518_U0_fifo_cout_drain_out_V_V_din,
  fifo_cout_drain_cout_drain_IO_L1_out_9_8_V_V_full_n,
  cout_drain_IO_L1_out_wrapper518_U0_fifo_cout_drain_out_V_V_write,
  PE_wrapper255_U0_fifo_cin_out_V_V_din,
  fifo_cin_PE_9_9_V_V_full_n,
  PE_wrapper255_U0_fifo_cin_out_V_V_write,
  PE_wrapper244_U0_fifo_w_out_V_V_din,
  fifo_w_PE_7_11_V_V_full_n,
  PE_wrapper244_U0_fifo_w_out_V_V_write,
  PE_wrapper173_U0_fifo_cout_drain_out_V_din,
  fifo_cout_drain_PE_1_11_V_full_n,
  PE_wrapper173_U0_fifo_cout_drain_out_V_write,
  PE_wrapper254_U0_fifo_w_out_V_V_din,
  fifo_w_PE_8_9_V_V_full_n,
  PE_wrapper254_U0_fifo_w_out_V_V_write,
  PE_wrapper208_U0_fifo_cout_drain_out_V_din,
  fifo_cout_drain_PE_4_10_V_full_n,
  PE_wrapper208_U0_fifo_cout_drain_out_V_write,
  cout_drain_IO_L1_out_wrapper536_U0_fifo_cout_drain_out_V_V_din,
  fifo_cout_drain_cout_drain_IO_L1_out_10_6_V_V_full_n,
  cout_drain_IO_L1_out_wrapper536_U0_fifo_cout_drain_out_V_V_write,
  PE_wrapper182_U0_fifo_w_out_V_V_din,
  fifo_w_PE_2_9_V_V_full_n,
  PE_wrapper182_U0_fifo_w_out_V_V_write,
  PE_wrapper220_U0_fifo_w_out_V_V_din,
  fifo_w_PE_5_11_V_V_full_n,
  PE_wrapper220_U0_fifo_w_out_V_V_write,
  PE_wrapper255_U0_fifo_w_out_V_V_din,
  fifo_w_PE_8_10_V_V_full_n,
  PE_wrapper255_U0_fifo_w_out_V_V_write,
  cout_drain_IO_L1_out_wrapper534_U0_fifo_cout_drain_out_V_V_din,
  fifo_cout_drain_cout_drain_IO_L1_out_10_8_V_V_full_n,
  cout_drain_IO_L1_out_wrapper534_U0_fifo_cout_drain_out_V_V_write,
  cout_drain_IO_L1_out_wrapper520_U0_fifo_cout_drain_out_V_V_din,
  fifo_cout_drain_cout_drain_IO_L1_out_9_6_V_V_full_n,
  cout_drain_IO_L1_out_wrapper520_U0_fifo_cout_drain_out_V_V_write,
  cout_drain_IO_L3_out_U0_fifo_cout_drain_out_V_V_din,
  fifo_cout_drain_cout_drain_IO_L3_out_serialize_V_V_full_n,
  cout_drain_IO_L3_out_U0_fifo_cout_drain_out_V_V_write,
  PE_wrapper173_U0_fifo_cin_out_V_V_din,
  fifo_cin_PE_2_11_V_V_full_n,
  PE_wrapper173_U0_fifo_cin_out_V_V_write,
  PE_wrapper232_U0_fifo_w_out_V_V_din,
  fifo_w_PE_6_11_V_V_full_n,
  PE_wrapper232_U0_fifo_w_out_V_V_write,
  PE_wrapper183_U0_fifo_w_out_V_V_din,
  fifo_w_PE_2_10_V_V_full_n,
  PE_wrapper183_U0_fifo_w_out_V_V_write,
  PE_wrapper221_U0_fifo_w_out_V_V_din,
  fifo_w_PE_5_12_V_V_full_n,
  PE_wrapper221_U0_fifo_w_out_V_V_write,
  PE_wrapper208_U0_fifo_w_out_V_V_din,
  fifo_w_PE_4_11_V_V_full_n,
  PE_wrapper208_U0_fifo_w_out_V_V_write,
  PE_wrapper197_U0_fifo_cout_drain_out_V_din,
  fifo_cout_drain_PE_3_11_V_full_n,
  PE_wrapper197_U0_fifo_cout_drain_out_V_write,
  PE_wrapper183_U0_fifo_cin_out_V_V_din,
  fifo_cin_PE_3_9_V_V_full_n,
  PE_wrapper183_U0_fifo_cin_out_V_V_write,
  cout_drain_IO_L1_out_wrapper553_U0_fifo_cout_drain_out_V_V_din,
  fifo_cout_drain_cout_drain_IO_L1_out_11_4_V_V_full_n,
  cout_drain_IO_L1_out_wrapper553_U0_fifo_cout_drain_out_V_V_write,
  m_axi_gmem_cout_AWVALID,
  m_axi_gmem_cout_AWREADY,
  m_axi_gmem_cout_AWADDR,
  m_axi_gmem_cout_AWID,
  m_axi_gmem_cout_AWLEN,
  m_axi_gmem_cout_AWSIZE,
  m_axi_gmem_cout_AWBURST,
  m_axi_gmem_cout_AWLOCK,
  m_axi_gmem_cout_AWCACHE,
  m_axi_gmem_cout_AWPROT,
  m_axi_gmem_cout_AWQOS,
  m_axi_gmem_cout_AWREGION,
  m_axi_gmem_cout_AWUSER,
  m_axi_gmem_cout_WVALID,
  m_axi_gmem_cout_WREADY,
  m_axi_gmem_cout_WDATA,
  m_axi_gmem_cout_WSTRB,
  m_axi_gmem_cout_WLAST,
  m_axi_gmem_cout_WID,
  m_axi_gmem_cout_WUSER,
  m_axi_gmem_cout_ARVALID,
  m_axi_gmem_cout_ARREADY,
  m_axi_gmem_cout_ARADDR,
  m_axi_gmem_cout_ARID,
  m_axi_gmem_cout_ARLEN,
  m_axi_gmem_cout_ARSIZE,
  m_axi_gmem_cout_ARBURST,
  m_axi_gmem_cout_ARLOCK,
  m_axi_gmem_cout_ARCACHE,
  m_axi_gmem_cout_ARPROT,
  m_axi_gmem_cout_ARQOS,
  m_axi_gmem_cout_ARREGION,
  m_axi_gmem_cout_ARUSER,
  m_axi_gmem_cout_RVALID,
  m_axi_gmem_cout_RREADY,
  m_axi_gmem_cout_RDATA,
  m_axi_gmem_cout_RLAST,
  m_axi_gmem_cout_RID,
  m_axi_gmem_cout_RUSER,
  m_axi_gmem_cout_RRESP,
  m_axi_gmem_cout_BVALID,
  m_axi_gmem_cout_BREADY,
  m_axi_gmem_cout_BRESP,
  m_axi_gmem_cout_BID,
  m_axi_gmem_cout_BUSER,
  ap_start,
  ap_done,
  ap_idle,
  ap_ready,
  ap_continue,
  ap_clk,
  ap_rst_n
);
parameter C_S_AXI_CONTROL_DATA_WIDTH = 32;
parameter C_S_AXI_CONTROL_ADDR_WIDTH = 6;
parameter C_S_AXI_DATA_WIDTH = 32;
parameter C_S_AXI_ADDR_WIDTH = 32;
parameter C_M_AXI_GMEM_CIN_ID_WIDTH = 1;
parameter C_M_AXI_GMEM_CIN_ADDR_WIDTH = 64;
parameter C_M_AXI_GMEM_CIN_DATA_WIDTH = 512;
parameter C_M_AXI_GMEM_CIN_AWUSER_WIDTH = 1;
parameter C_M_AXI_GMEM_CIN_ARUSER_WIDTH = 1;
parameter C_M_AXI_GMEM_CIN_WUSER_WIDTH = 1;
parameter C_M_AXI_GMEM_CIN_RUSER_WIDTH = 1;
parameter C_M_AXI_GMEM_CIN_BUSER_WIDTH = 1;
parameter C_M_AXI_GMEM_CIN_USER_VALUE = 0;
parameter C_M_AXI_GMEM_CIN_PROT_VALUE = 0;
parameter C_M_AXI_GMEM_CIN_CACHE_VALUE = 3;
parameter C_M_AXI_ID_WIDTH = 1;
parameter C_M_AXI_ADDR_WIDTH = 64;
parameter C_M_AXI_DATA_WIDTH = 32;
parameter C_M_AXI_AWUSER_WIDTH = 1;
parameter C_M_AXI_ARUSER_WIDTH = 1;
parameter C_M_AXI_WUSER_WIDTH = 1;
parameter C_M_AXI_RUSER_WIDTH = 1;
parameter C_M_AXI_BUSER_WIDTH = 1;
parameter C_M_AXI_GMEM_COUT_ID_WIDTH = 1;
parameter C_M_AXI_GMEM_COUT_ADDR_WIDTH = 64;
parameter C_M_AXI_GMEM_COUT_DATA_WIDTH = 512;
parameter C_M_AXI_GMEM_COUT_AWUSER_WIDTH = 1;
parameter C_M_AXI_GMEM_COUT_ARUSER_WIDTH = 1;
parameter C_M_AXI_GMEM_COUT_WUSER_WIDTH = 1;
parameter C_M_AXI_GMEM_COUT_RUSER_WIDTH = 1;
parameter C_M_AXI_GMEM_COUT_BUSER_WIDTH = 1;
parameter C_M_AXI_GMEM_COUT_USER_VALUE = 0;
parameter C_M_AXI_GMEM_COUT_PROT_VALUE = 0;
parameter C_M_AXI_GMEM_COUT_CACHE_VALUE = 3;
parameter C_M_AXI_GMEM_W_ID_WIDTH = 1;
parameter C_M_AXI_GMEM_W_ADDR_WIDTH = 64;
parameter C_M_AXI_GMEM_W_DATA_WIDTH = 512;
parameter C_M_AXI_GMEM_W_AWUSER_WIDTH = 1;
parameter C_M_AXI_GMEM_W_ARUSER_WIDTH = 1;
parameter C_M_AXI_GMEM_W_WUSER_WIDTH = 1;
parameter C_M_AXI_GMEM_W_RUSER_WIDTH = 1;
parameter C_M_AXI_GMEM_W_BUSER_WIDTH = 1;
parameter C_M_AXI_GMEM_W_USER_VALUE = 0;
parameter C_M_AXI_GMEM_W_PROT_VALUE = 0;
parameter C_M_AXI_GMEM_W_CACHE_VALUE = 3;
parameter C_S_AXI_CONTROL_WSTRB_WIDTH = 32 / 8;
parameter C_S_AXI_WSTRB_WIDTH = 32 / 8;
parameter C_M_AXI_GMEM_CIN_WSTRB_WIDTH = 512 / 8;
parameter C_M_AXI_WSTRB_WIDTH = 32 / 8;
parameter C_M_AXI_GMEM_COUT_WSTRB_WIDTH = 512 / 8;
parameter C_M_AXI_GMEM_W_WSTRB_WIDTH = 512 / 8;
reg ap_rst_n_inv;
wire gmem_cout_AWREADY;
wire gmem_cout_WREADY;
wire gmem_cout_ARREADY;
wire gmem_cout_RVALID;
wire [511:0] gmem_cout_RDATA;
wire gmem_cout_RLAST;
wire [0:0] gmem_cout_RID;
wire [0:0] gmem_cout_RUSER;
wire [1:0] gmem_cout_RRESP;
wire gmem_cout_BVALID;
wire [1:0] gmem_cout_BRESP;
wire [0:0] gmem_cout_BID;
wire [0:0] gmem_cout_BUSER;
wire PE_wrapper173_U0_ap_start;
wire PE_wrapper173_U0_ap_done;
wire PE_wrapper173_U0_ap_continue;
wire PE_wrapper173_U0_ap_idle;
wire PE_wrapper173_U0_ap_ready;
wire PE_wrapper173_U0_fifo_cin_in_V_V_read;
wire PE_wrapper173_U0_fifo_w_in_V_V_read;
wire PE_wrapper183_U0_ap_start;
wire PE_wrapper183_U0_ap_done;
wire PE_wrapper183_U0_ap_continue;
wire PE_wrapper183_U0_ap_idle;
wire PE_wrapper183_U0_ap_ready;
wire PE_wrapper183_U0_fifo_cin_in_V_V_read;
wire PE_wrapper183_U0_fifo_w_in_V_V_read;
wire PE_wrapper208_U0_ap_start;
wire PE_wrapper208_U0_ap_done;
wire PE_wrapper208_U0_ap_continue;
wire PE_wrapper208_U0_ap_idle;
wire PE_wrapper208_U0_ap_ready;
wire PE_wrapper208_U0_fifo_cin_in_V_V_read;
wire [255:0] PE_wrapper208_U0_fifo_cin_out_V_V_din;
wire PE_wrapper208_U0_fifo_cin_out_V_V_write;
wire PE_wrapper208_U0_fifo_w_in_V_V_read;
wire PE_wrapper220_U0_ap_start;
wire PE_wrapper220_U0_ap_done;
wire PE_wrapper220_U0_ap_continue;
wire PE_wrapper220_U0_ap_idle;
wire PE_wrapper220_U0_ap_ready;
wire PE_wrapper220_U0_fifo_cin_in_V_V_read;
wire [255:0] PE_wrapper220_U0_fifo_cin_out_V_V_din;
wire PE_wrapper220_U0_fifo_cin_out_V_V_write;
wire [31:0] PE_wrapper220_U0_fifo_cout_drain_out_V_din;
wire PE_wrapper220_U0_fifo_cout_drain_out_V_write;
wire PE_wrapper220_U0_fifo_w_in_V_V_read;
wire PE_wrapper232_U0_ap_start;
wire PE_wrapper232_U0_ap_done;
wire PE_wrapper232_U0_ap_continue;
wire PE_wrapper232_U0_ap_idle;
wire PE_wrapper232_U0_ap_ready;
wire PE_wrapper232_U0_fifo_cin_in_V_V_read;
wire [255:0] PE_wrapper232_U0_fifo_cin_out_V_V_din;
wire PE_wrapper232_U0_fifo_cin_out_V_V_write;
wire PE_wrapper232_U0_fifo_w_in_V_V_read;
wire PE_wrapper244_U0_ap_start;
wire PE_wrapper244_U0_ap_done;
wire PE_wrapper244_U0_ap_continue;
wire PE_wrapper244_U0_ap_idle;
wire PE_wrapper244_U0_ap_ready;
wire PE_wrapper244_U0_fifo_cin_in_V_V_read;
wire [31:0] PE_wrapper244_U0_fifo_cout_drain_out_V_din;
wire PE_wrapper244_U0_fifo_cout_drain_out_V_write;
wire PE_wrapper244_U0_fifo_w_in_V_V_read;
wire PE_wrapper255_U0_ap_start;
wire PE_wrapper255_U0_ap_done;
wire PE_wrapper255_U0_ap_continue;
wire PE_wrapper255_U0_ap_idle;
wire PE_wrapper255_U0_ap_ready;
wire PE_wrapper255_U0_fifo_cin_in_V_V_read;
wire PE_wrapper255_U0_fifo_w_in_V_V_read;
wire w_PE_dummy_in357_U0_ap_start;
wire w_PE_dummy_in357_U0_ap_done;
wire w_PE_dummy_in357_U0_ap_continue;
wire w_PE_dummy_in357_U0_ap_idle;
wire w_PE_dummy_in357_U0_ap_ready;
wire w_PE_dummy_in357_U0_fifo_w_in_V_V_read;
wire cout_drain_IO_L1_out_wrapper519_U0_ap_start;
wire cout_drain_IO_L1_out_wrapper519_U0_ap_done;
wire cout_drain_IO_L1_out_wrapper519_U0_ap_continue;
wire cout_drain_IO_L1_out_wrapper519_U0_ap_idle;
wire cout_drain_IO_L1_out_wrapper519_U0_ap_ready;
wire cout_drain_IO_L1_out_wrapper519_U0_fifo_cout_drain_in_V_V_read;
wire [63:0] cout_drain_IO_L1_out_wrapper519_U0_fifo_cout_drain_out_V_V_din;
wire cout_drain_IO_L1_out_wrapper519_U0_fifo_cout_drain_out_V_V_write;
wire cout_drain_IO_L1_out_wrapper519_U0_fifo_cout_drain_local_in_V_read;
wire cout_drain_IO_L1_out_wrapper520_U0_ap_start;
wire cout_drain_IO_L1_out_wrapper520_U0_ap_done;
wire cout_drain_IO_L1_out_wrapper520_U0_ap_continue;
wire cout_drain_IO_L1_out_wrapper520_U0_ap_idle;
wire cout_drain_IO_L1_out_wrapper520_U0_ap_ready;
wire cout_drain_IO_L1_out_wrapper520_U0_fifo_cout_drain_in_V_V_read;
wire cout_drain_IO_L1_out_wrapper520_U0_fifo_cout_drain_local_in_V_read;
wire cout_drain_IO_L1_out_wrapper535_U0_ap_start;
wire cout_drain_IO_L1_out_wrapper535_U0_ap_done;
wire cout_drain_IO_L1_out_wrapper535_U0_ap_continue;
wire cout_drain_IO_L1_out_wrapper535_U0_ap_idle;
wire cout_drain_IO_L1_out_wrapper535_U0_ap_ready;
wire cout_drain_IO_L1_out_wrapper535_U0_fifo_cout_drain_in_V_V_read;
wire cout_drain_IO_L1_out_wrapper535_U0_fifo_cout_drain_local_in_V_read;
wire cout_drain_IO_L1_out_wrapper537_U0_ap_start;
wire cout_drain_IO_L1_out_wrapper537_U0_ap_done;
wire cout_drain_IO_L1_out_wrapper537_U0_ap_continue;
wire cout_drain_IO_L1_out_wrapper537_U0_ap_idle;
wire cout_drain_IO_L1_out_wrapper537_U0_ap_ready;
wire cout_drain_IO_L1_out_wrapper537_U0_fifo_cout_drain_in_V_V_read;
wire cout_drain_IO_L1_out_wrapper537_U0_fifo_cout_drain_local_in_V_read;
wire cout_drain_IO_L1_out_wrapper540_U0_ap_start;
wire cout_drain_IO_L1_out_wrapper540_U0_ap_done;
wire cout_drain_IO_L1_out_wrapper540_U0_ap_continue;
wire cout_drain_IO_L1_out_wrapper540_U0_ap_idle;
wire cout_drain_IO_L1_out_wrapper540_U0_ap_ready;
wire cout_drain_IO_L1_out_wrapper540_U0_fifo_cout_drain_in_V_V_read;
wire cout_drain_IO_L1_out_wrapper540_U0_fifo_cout_drain_local_in_V_read;
wire cout_drain_IO_L1_out_wrapper552_U0_ap_start;
wire cout_drain_IO_L1_out_wrapper552_U0_ap_done;
wire cout_drain_IO_L1_out_wrapper552_U0_ap_continue;
wire cout_drain_IO_L1_out_wrapper552_U0_ap_idle;
wire cout_drain_IO_L1_out_wrapper552_U0_ap_ready;
wire cout_drain_IO_L1_out_wrapper552_U0_fifo_cout_drain_in_V_V_read;
wire cout_drain_IO_L1_out_wrapper552_U0_fifo_cout_drain_local_in_V_read;
wire cout_drain_IO_L1_out_wrapper554_U0_ap_start;
wire cout_drain_IO_L1_out_wrapper554_U0_ap_done;
wire cout_drain_IO_L1_out_wrapper554_U0_ap_continue;
wire cout_drain_IO_L1_out_wrapper554_U0_ap_idle;
wire cout_drain_IO_L1_out_wrapper554_U0_ap_ready;
wire cout_drain_IO_L1_out_wrapper554_U0_fifo_cout_drain_in_V_V_read;
wire [63:0] cout_drain_IO_L1_out_wrapper554_U0_fifo_cout_drain_out_V_V_din;
wire cout_drain_IO_L1_out_wrapper554_U0_fifo_cout_drain_out_V_V_write;
wire cout_drain_IO_L1_out_wrapper554_U0_fifo_cout_drain_local_in_V_read;
wire cout_drain_IO_L1_out_wrapper555_U0_ap_start;
wire cout_drain_IO_L1_out_wrapper555_U0_ap_done;
wire cout_drain_IO_L1_out_wrapper555_U0_ap_continue;
wire cout_drain_IO_L1_out_wrapper555_U0_ap_idle;
wire cout_drain_IO_L1_out_wrapper555_U0_ap_ready;
wire cout_drain_IO_L1_out_wrapper555_U0_fifo_cout_drain_in_V_V_read;
wire cout_drain_IO_L1_out_wrapper555_U0_fifo_cout_drain_local_in_V_read;
wire cout_drain_IO_L3_out_serialize_U0_ap_start;
wire cout_drain_IO_L3_out_serialize_U0_ap_done;
wire cout_drain_IO_L3_out_serialize_U0_ap_continue;
wire cout_drain_IO_L3_out_serialize_U0_ap_idle;
wire cout_drain_IO_L3_out_serialize_U0_ap_ready;
wire cout_drain_IO_L3_out_serialize_U0_m_axi_cout_V_AWVALID;
wire [63:0] cout_drain_IO_L3_out_serialize_U0_m_axi_cout_V_AWADDR;
wire [0:0] cout_drain_IO_L3_out_serialize_U0_m_axi_cout_V_AWID;
wire [31:0] cout_drain_IO_L3_out_serialize_U0_m_axi_cout_V_AWLEN;
wire [2:0] cout_drain_IO_L3_out_serialize_U0_m_axi_cout_V_AWSIZE;
wire [1:0] cout_drain_IO_L3_out_serialize_U0_m_axi_cout_V_AWBURST;
wire [1:0] cout_drain_IO_L3_out_serialize_U0_m_axi_cout_V_AWLOCK;
wire [3:0] cout_drain_IO_L3_out_serialize_U0_m_axi_cout_V_AWCACHE;
wire [2:0] cout_drain_IO_L3_out_serialize_U0_m_axi_cout_V_AWPROT;
wire [3:0] cout_drain_IO_L3_out_serialize_U0_m_axi_cout_V_AWQOS;
wire [3:0] cout_drain_IO_L3_out_serialize_U0_m_axi_cout_V_AWREGION;
wire [0:0] cout_drain_IO_L3_out_serialize_U0_m_axi_cout_V_AWUSER;
wire cout_drain_IO_L3_out_serialize_U0_m_axi_cout_V_WVALID;
wire [511:0] cout_drain_IO_L3_out_serialize_U0_m_axi_cout_V_WDATA;
wire [63:0] cout_drain_IO_L3_out_serialize_U0_m_axi_cout_V_WSTRB;
wire cout_drain_IO_L3_out_serialize_U0_m_axi_cout_V_WLAST;
wire [0:0] cout_drain_IO_L3_out_serialize_U0_m_axi_cout_V_WID;
wire [0:0] cout_drain_IO_L3_out_serialize_U0_m_axi_cout_V_WUSER;
wire cout_drain_IO_L3_out_serialize_U0_m_axi_cout_V_ARVALID;
wire [63:0] cout_drain_IO_L3_out_serialize_U0_m_axi_cout_V_ARADDR;
wire [0:0] cout_drain_IO_L3_out_serialize_U0_m_axi_cout_V_ARID;
wire [31:0] cout_drain_IO_L3_out_serialize_U0_m_axi_cout_V_ARLEN;
wire [2:0] cout_drain_IO_L3_out_serialize_U0_m_axi_cout_V_ARSIZE;
wire [1:0] cout_drain_IO_L3_out_serialize_U0_m_axi_cout_V_ARBURST;
wire [1:0] cout_drain_IO_L3_out_serialize_U0_m_axi_cout_V_ARLOCK;
wire [3:0] cout_drain_IO_L3_out_serialize_U0_m_axi_cout_V_ARCACHE;
wire [2:0] cout_drain_IO_L3_out_serialize_U0_m_axi_cout_V_ARPROT;
wire [3:0] cout_drain_IO_L3_out_serialize_U0_m_axi_cout_V_ARQOS;
wire [3:0] cout_drain_IO_L3_out_serialize_U0_m_axi_cout_V_ARREGION;
wire [0:0] cout_drain_IO_L3_out_serialize_U0_m_axi_cout_V_ARUSER;
wire cout_drain_IO_L3_out_serialize_U0_m_axi_cout_V_RREADY;
wire cout_drain_IO_L3_out_serialize_U0_m_axi_cout_V_BREADY;
wire cout_drain_IO_L3_out_serialize_U0_cout_V_offset_read;
wire cout_drain_IO_L3_out_serialize_U0_fifo_cout_drain_local_in_V_V_read;
wire [63:0] cout_V_c_dout;
wire cout_V_c_empty_n;
wire [255:0] fifo_cin_PE_1_11_V_V_dout;
wire fifo_cin_PE_1_11_V_V_empty_n;
wire [255:0] fifo_cin_PE_2_9_V_V_dout;
wire fifo_cin_PE_2_9_V_V_empty_n;
wire [255:0] fifo_w_PE_1_11_V_V_dout;
wire fifo_w_PE_1_11_V_V_empty_n;
wire [255:0] fifo_w_PE_2_9_V_V_dout;
wire fifo_w_PE_2_9_V_V_empty_n;
wire [31:0] fifo_cout_drain_PE_2_10_V_dout;
wire fifo_cout_drain_PE_2_10_V_empty_n;
wire [31:0] fifo_cout_drain_PE_2_11_V_dout;
wire fifo_cout_drain_PE_2_11_V_empty_n;
wire [255:0] fifo_cin_PE_4_10_V_V_dout;
wire fifo_cin_PE_4_10_V_V_empty_n;
wire [31:0] fifo_cout_drain_PE_3_11_V_dout;
wire fifo_cout_drain_PE_3_11_V_empty_n;
wire [255:0] fifo_w_PE_4_10_V_V_dout;
wire fifo_w_PE_4_10_V_V_empty_n;
wire fifo_cin_PE_5_10_V_V_full_n;
wire [255:0] fifo_cin_PE_5_10_V_V_dout;
wire fifo_cin_PE_5_10_V_V_empty_n;
wire [255:0] fifo_w_PE_5_10_V_V_dout;
wire fifo_w_PE_5_10_V_V_empty_n;
wire fifo_cin_PE_6_10_V_V_full_n;
wire [255:0] fifo_cin_PE_6_10_V_V_dout;
wire fifo_cin_PE_6_10_V_V_empty_n;
wire fifo_cout_drain_PE_5_10_V_full_n;
wire [31:0] fifo_cout_drain_PE_5_10_V_dout;
wire fifo_cout_drain_PE_5_10_V_empty_n;
wire [31:0] fifo_cout_drain_PE_5_11_V_dout;
wire fifo_cout_drain_PE_5_11_V_empty_n;
wire [255:0] fifo_w_PE_5_12_V_V_dout;
wire fifo_w_PE_5_12_V_V_empty_n;
wire [31:0] fifo_cout_drain_PE_6_9_V_dout;
wire fifo_cout_drain_PE_6_9_V_empty_n;
wire [255:0] fifo_w_PE_6_10_V_V_dout;
wire fifo_w_PE_6_10_V_V_empty_n;
wire fifo_cin_PE_7_10_V_V_full_n;
wire [255:0] fifo_cin_PE_7_10_V_V_dout;
wire fifo_cin_PE_7_10_V_V_empty_n;
wire [255:0] fifo_cin_PE_8_9_V_V_dout;
wire fifo_cin_PE_8_9_V_V_empty_n;
wire [31:0] fifo_cout_drain_PE_7_9_V_dout;
wire fifo_cout_drain_PE_7_9_V_empty_n;
wire [255:0] fifo_w_PE_7_10_V_V_dout;
wire fifo_w_PE_7_10_V_V_empty_n;
wire fifo_cout_drain_PE_7_10_V_full_n;
wire [31:0] fifo_cout_drain_PE_7_10_V_dout;
wire fifo_cout_drain_PE_7_10_V_empty_n;
wire [255:0] fifo_w_PE_8_9_V_V_dout;
wire fifo_w_PE_8_9_V_V_empty_n;
wire [63:0] fifo_cout_drain_cout_drain_IO_L1_out_9_8_V_V_dout;
wire fifo_cout_drain_cout_drain_IO_L1_out_9_8_V_V_empty_n;
wire fifo_cout_drain_cout_drain_IO_L1_out_9_7_V_V_full_n;
wire [63:0] fifo_cout_drain_cout_drain_IO_L1_out_9_7_V_V_dout;
wire fifo_cout_drain_cout_drain_IO_L1_out_9_7_V_V_empty_n;
wire [63:0] fifo_cout_drain_cout_drain_IO_L1_out_10_8_V_V_dout;
wire fifo_cout_drain_cout_drain_IO_L1_out_10_8_V_V_empty_n;
wire [63:0] fifo_cout_drain_cout_drain_IO_L1_out_10_6_V_V_dout;
wire fifo_cout_drain_cout_drain_IO_L1_out_10_6_V_V_empty_n;
wire [63:0] fifo_cout_drain_cout_drain_IO_L1_out_10_3_V_V_dout;
wire fifo_cout_drain_cout_drain_IO_L1_out_10_3_V_V_empty_n;
wire [63:0] fifo_cout_drain_cout_drain_IO_L1_out_11_6_V_V_dout;
wire fifo_cout_drain_cout_drain_IO_L1_out_11_6_V_V_empty_n;
wire [63:0] fifo_cout_drain_cout_drain_IO_L1_out_11_4_V_V_dout;
wire fifo_cout_drain_cout_drain_IO_L1_out_11_4_V_V_empty_n;
wire fifo_cout_drain_cout_drain_IO_L1_out_11_3_V_V_full_n;
wire [63:0] fifo_cout_drain_cout_drain_IO_L1_out_11_3_V_V_dout;
wire fifo_cout_drain_cout_drain_IO_L1_out_11_3_V_V_empty_n;
wire [63:0] fifo_cout_drain_cout_drain_IO_L3_out_serialize_V_V_dout;
wire fifo_cout_drain_cout_drain_IO_L3_out_serialize_V_V_empty_n;
// pipeline ap_start
(* shreg_extract = "no" *) reg ap_start_p1;
(* shreg_extract = "no" *) reg ap_start_p2;
(* shreg_extract = "no" *) reg ap_start_pipe;
// pipeline ap_done
(* shreg_extract = "no" *) reg w_PE_dummy_in357_U0_ap_done_p1;
(* shreg_extract = "no" *) reg w_PE_dummy_in357_U0_ap_done_p2;
(* shreg_extract = "no" *) reg w_PE_dummy_in357_U0_ap_done_pipe;
(* shreg_extract = "no" *) reg w_PE_dummy_in357_U0_ap_done_backup;
(* shreg_extract = "no" *) reg cout_drain_IO_L3_out_serialize_U0_ap_done_p1;
(* shreg_extract = "no" *) reg cout_drain_IO_L3_out_serialize_U0_ap_done_p2;
(* shreg_extract = "no" *) reg cout_drain_IO_L3_out_serialize_U0_ap_done_pipe;
(* shreg_extract = "no" *) reg cout_drain_IO_L3_out_serialize_U0_ap_done_backup;
// pipeline ap_rst_n
(* shreg_extract = "no" *) reg ap_rst_p1;
(* shreg_extract = "no" *) reg ap_rst_p2;
(* shreg_extract = "no" *) reg ap_rst_pipe;
(* shreg_extract = "no" *) reg ap_rst_n_p1;
(* shreg_extract = "no" *) reg ap_rst_n_p2;
(* shreg_extract = "no" *) reg ap_rst_n_pipe;
output [63:0] cout_drain_IO_L1_out_wrapper535_U0_fifo_cout_drain_out_V_V_din;
input  fifo_cout_drain_cout_drain_IO_L1_out_10_7_V_V_full_n;
output  cout_drain_IO_L1_out_wrapper535_U0_fifo_cout_drain_out_V_V_write;
input [255:0] PE_wrapper219_U0_fifo_w_out_V_V_din;
output  fifo_w_PE_5_10_V_V_full_n;
input  PE_wrapper219_U0_fifo_w_out_V_V_write;
output [63:0] cout_drain_IO_L1_out_wrapper537_U0_fifo_cout_drain_out_V_V_din;
input  fifo_cout_drain_cout_drain_IO_L1_out_10_5_V_V_full_n;
output  cout_drain_IO_L1_out_wrapper537_U0_fifo_cout_drain_out_V_V_write;
input [255:0] PE_wrapper171_U0_fifo_cin_out_V_V_din;
output  fifo_cin_PE_2_9_V_V_full_n;
input  PE_wrapper171_U0_fifo_cin_out_V_V_write;
input [255:0] PE_wrapper172_U0_fifo_w_out_V_V_din;
output  fifo_w_PE_1_11_V_V_full_n;
input  PE_wrapper172_U0_fifo_w_out_V_V_write;
input [63:0] cout_drain_IO_L1_out_wrapper551_U0_fifo_cout_drain_out_V_V_din;
output  fifo_cout_drain_cout_drain_IO_L1_out_11_6_V_V_full_n;
input  cout_drain_IO_L1_out_wrapper551_U0_fifo_cout_drain_out_V_V_write;
output [63:0] cout_drain_IO_L1_out_wrapper555_U0_fifo_cout_drain_out_V_V_din;
input  fifo_cout_drain_cout_drain_IO_L1_out_11_2_V_V_full_n;
output  cout_drain_IO_L1_out_wrapper555_U0_fifo_cout_drain_out_V_V_write;
input [255:0] PE_wrapper196_U0_fifo_cin_out_V_V_din;
output  fifo_cin_PE_4_10_V_V_full_n;
input  PE_wrapper196_U0_fifo_cin_out_V_V_write;
input [63:0] cout_drain_IO_L1_out_wrapper539_U0_fifo_cout_drain_out_V_V_din;
output  fifo_cout_drain_cout_drain_IO_L1_out_10_3_V_V_full_n;
input  cout_drain_IO_L1_out_wrapper539_U0_fifo_cout_drain_out_V_V_write;
output [255:0] PE_wrapper244_U0_fifo_cin_out_V_V_din;
input  fifo_cin_PE_8_10_V_V_full_n;
output  PE_wrapper244_U0_fifo_cin_out_V_V_write;
input [255:0] PE_wrapper231_U0_fifo_w_out_V_V_din;
output  fifo_w_PE_6_10_V_V_full_n;
input  PE_wrapper231_U0_fifo_w_out_V_V_write;
output [255:0] PE_wrapper173_U0_fifo_w_out_V_V_din;
input  fifo_w_PE_1_12_V_V_full_n;
output  PE_wrapper173_U0_fifo_w_out_V_V_write;
input [31:0] PE_wrapper231_U0_fifo_cout_drain_out_V_din;
output  fifo_cout_drain_PE_6_9_V_full_n;
input  PE_wrapper231_U0_fifo_cout_drain_out_V_write;
input [255:0] PE_wrapper207_U0_fifo_w_out_V_V_din;
output  fifo_w_PE_4_10_V_V_full_n;
input  PE_wrapper207_U0_fifo_w_out_V_V_write;
input [31:0] PE_wrapper221_U0_fifo_cout_drain_out_V_din;
output  fifo_cout_drain_PE_5_11_V_full_n;
input  PE_wrapper221_U0_fifo_cout_drain_out_V_write;
output [31:0] PE_wrapper183_U0_fifo_cout_drain_out_V_din;
input  fifo_cout_drain_PE_2_9_V_full_n;
output  PE_wrapper183_U0_fifo_cout_drain_out_V_write;
input [255:0] PE_wrapper161_U0_fifo_cin_out_V_V_din;
output  fifo_cin_PE_1_11_V_V_full_n;
input  PE_wrapper161_U0_fifo_cin_out_V_V_write;
output [31:0] PE_wrapper232_U0_fifo_cout_drain_out_V_din;
input  fifo_cout_drain_PE_6_10_V_full_n;
output  PE_wrapper232_U0_fifo_cout_drain_out_V_write;
input [63:0] kernel0_entry12_U0_cout_V_out_din;
output  cout_V_c_full_n;
input  kernel0_entry12_U0_cout_V_out_write;
output [63:0] cout_drain_IO_L1_out_wrapper540_U0_fifo_cout_drain_out_V_V_din;
input  fifo_cout_drain_cout_drain_IO_L1_out_10_2_V_V_full_n;
output  cout_drain_IO_L1_out_wrapper540_U0_fifo_cout_drain_out_V_V_write;
output [63:0] cout_drain_IO_L1_out_wrapper552_U0_fifo_cout_drain_out_V_V_din;
input  fifo_cout_drain_cout_drain_IO_L1_out_11_5_V_V_full_n;
output  cout_drain_IO_L1_out_wrapper552_U0_fifo_cout_drain_out_V_V_write;
input [255:0] PE_wrapper243_U0_fifo_w_out_V_V_din;
output  fifo_w_PE_7_10_V_V_full_n;
input  PE_wrapper243_U0_fifo_w_out_V_V_write;
input [31:0] PE_wrapper243_U0_fifo_cout_drain_out_V_din;
output  fifo_cout_drain_PE_7_9_V_full_n;
input  PE_wrapper243_U0_fifo_cout_drain_out_V_write;
input [31:0] PE_wrapper184_U0_fifo_cout_drain_out_V_din;
output  fifo_cout_drain_PE_2_10_V_full_n;
input  PE_wrapper184_U0_fifo_cout_drain_out_V_write;
input [255:0] PE_wrapper243_U0_fifo_cin_out_V_V_din;
output  fifo_cin_PE_8_9_V_V_full_n;
input  PE_wrapper243_U0_fifo_cin_out_V_V_write;
output [31:0] PE_wrapper255_U0_fifo_cout_drain_out_V_din;
input  fifo_cout_drain_PE_8_9_V_full_n;
output  PE_wrapper255_U0_fifo_cout_drain_out_V_write;
input [31:0] PE_wrapper185_U0_fifo_cout_drain_out_V_din;
output  fifo_cout_drain_PE_2_11_V_full_n;
input  PE_wrapper185_U0_fifo_cout_drain_out_V_write;
input [63:0] cout_drain_IO_L1_out_wrapper518_U0_fifo_cout_drain_out_V_V_din;
output  fifo_cout_drain_cout_drain_IO_L1_out_9_8_V_V_full_n;
input  cout_drain_IO_L1_out_wrapper518_U0_fifo_cout_drain_out_V_V_write;
output [255:0] PE_wrapper255_U0_fifo_cin_out_V_V_din;
input  fifo_cin_PE_9_9_V_V_full_n;
output  PE_wrapper255_U0_fifo_cin_out_V_V_write;
output [255:0] PE_wrapper244_U0_fifo_w_out_V_V_din;
input  fifo_w_PE_7_11_V_V_full_n;
output  PE_wrapper244_U0_fifo_w_out_V_V_write;
output [31:0] PE_wrapper173_U0_fifo_cout_drain_out_V_din;
input  fifo_cout_drain_PE_1_11_V_full_n;
output  PE_wrapper173_U0_fifo_cout_drain_out_V_write;
input [255:0] PE_wrapper254_U0_fifo_w_out_V_V_din;
output  fifo_w_PE_8_9_V_V_full_n;
input  PE_wrapper254_U0_fifo_w_out_V_V_write;
output [31:0] PE_wrapper208_U0_fifo_cout_drain_out_V_din;
input  fifo_cout_drain_PE_4_10_V_full_n;
output  PE_wrapper208_U0_fifo_cout_drain_out_V_write;
input [63:0] cout_drain_IO_L1_out_wrapper536_U0_fifo_cout_drain_out_V_V_din;
output  fifo_cout_drain_cout_drain_IO_L1_out_10_6_V_V_full_n;
input  cout_drain_IO_L1_out_wrapper536_U0_fifo_cout_drain_out_V_V_write;
input [255:0] PE_wrapper182_U0_fifo_w_out_V_V_din;
output  fifo_w_PE_2_9_V_V_full_n;
input  PE_wrapper182_U0_fifo_w_out_V_V_write;
output [255:0] PE_wrapper220_U0_fifo_w_out_V_V_din;
input  fifo_w_PE_5_11_V_V_full_n;
output  PE_wrapper220_U0_fifo_w_out_V_V_write;
output [255:0] PE_wrapper255_U0_fifo_w_out_V_V_din;
input  fifo_w_PE_8_10_V_V_full_n;
output  PE_wrapper255_U0_fifo_w_out_V_V_write;
input [63:0] cout_drain_IO_L1_out_wrapper534_U0_fifo_cout_drain_out_V_V_din;
output  fifo_cout_drain_cout_drain_IO_L1_out_10_8_V_V_full_n;
input  cout_drain_IO_L1_out_wrapper534_U0_fifo_cout_drain_out_V_V_write;
output [63:0] cout_drain_IO_L1_out_wrapper520_U0_fifo_cout_drain_out_V_V_din;
input  fifo_cout_drain_cout_drain_IO_L1_out_9_6_V_V_full_n;
output  cout_drain_IO_L1_out_wrapper520_U0_fifo_cout_drain_out_V_V_write;
input [63:0] cout_drain_IO_L3_out_U0_fifo_cout_drain_out_V_V_din;
output  fifo_cout_drain_cout_drain_IO_L3_out_serialize_V_V_full_n;
input  cout_drain_IO_L3_out_U0_fifo_cout_drain_out_V_V_write;
output [255:0] PE_wrapper173_U0_fifo_cin_out_V_V_din;
input  fifo_cin_PE_2_11_V_V_full_n;
output  PE_wrapper173_U0_fifo_cin_out_V_V_write;
output [255:0] PE_wrapper232_U0_fifo_w_out_V_V_din;
input  fifo_w_PE_6_11_V_V_full_n;
output  PE_wrapper232_U0_fifo_w_out_V_V_write;
output [255:0] PE_wrapper183_U0_fifo_w_out_V_V_din;
input  fifo_w_PE_2_10_V_V_full_n;
output  PE_wrapper183_U0_fifo_w_out_V_V_write;
input [255:0] PE_wrapper221_U0_fifo_w_out_V_V_din;
output  fifo_w_PE_5_12_V_V_full_n;
input  PE_wrapper221_U0_fifo_w_out_V_V_write;
output [255:0] PE_wrapper208_U0_fifo_w_out_V_V_din;
input  fifo_w_PE_4_11_V_V_full_n;
output  PE_wrapper208_U0_fifo_w_out_V_V_write;
input [31:0] PE_wrapper197_U0_fifo_cout_drain_out_V_din;
output  fifo_cout_drain_PE_3_11_V_full_n;
input  PE_wrapper197_U0_fifo_cout_drain_out_V_write;
output [255:0] PE_wrapper183_U0_fifo_cin_out_V_V_din;
input  fifo_cin_PE_3_9_V_V_full_n;
output  PE_wrapper183_U0_fifo_cin_out_V_V_write;
input [63:0] cout_drain_IO_L1_out_wrapper553_U0_fifo_cout_drain_out_V_V_din;
output  fifo_cout_drain_cout_drain_IO_L1_out_11_4_V_V_full_n;
input  cout_drain_IO_L1_out_wrapper553_U0_fifo_cout_drain_out_V_V_write;
output  m_axi_gmem_cout_AWVALID;
input  m_axi_gmem_cout_AWREADY;
output [64-1:0] m_axi_gmem_cout_AWADDR;
output [1-1:0] m_axi_gmem_cout_AWID;
output [7:0] m_axi_gmem_cout_AWLEN;
output [2:0] m_axi_gmem_cout_AWSIZE;
output [1:0] m_axi_gmem_cout_AWBURST;
output [1:0] m_axi_gmem_cout_AWLOCK;
output [3:0] m_axi_gmem_cout_AWCACHE;
output [2:0] m_axi_gmem_cout_AWPROT;
output [3:0] m_axi_gmem_cout_AWQOS;
output [3:0] m_axi_gmem_cout_AWREGION;
output [1-1:0] m_axi_gmem_cout_AWUSER;
output  m_axi_gmem_cout_WVALID;
input  m_axi_gmem_cout_WREADY;
output [512-1:0] m_axi_gmem_cout_WDATA;
output [512/8-1:0] m_axi_gmem_cout_WSTRB;
output  m_axi_gmem_cout_WLAST;
output [1-1:0] m_axi_gmem_cout_WID;
output [1-1:0] m_axi_gmem_cout_WUSER;
output  m_axi_gmem_cout_ARVALID;
input  m_axi_gmem_cout_ARREADY;
output [64-1:0] m_axi_gmem_cout_ARADDR;
output [1-1:0] m_axi_gmem_cout_ARID;
output [7:0] m_axi_gmem_cout_ARLEN;
output [2:0] m_axi_gmem_cout_ARSIZE;
output [1:0] m_axi_gmem_cout_ARBURST;
output [1:0] m_axi_gmem_cout_ARLOCK;
output [3:0] m_axi_gmem_cout_ARCACHE;
output [2:0] m_axi_gmem_cout_ARPROT;
output [3:0] m_axi_gmem_cout_ARQOS;
output [3:0] m_axi_gmem_cout_ARREGION;
output [1-1:0] m_axi_gmem_cout_ARUSER;
input  m_axi_gmem_cout_RVALID;
output  m_axi_gmem_cout_RREADY;
input [512-1:0] m_axi_gmem_cout_RDATA;
input  m_axi_gmem_cout_RLAST;
input [1-1:0] m_axi_gmem_cout_RID;
input [1-1:0] m_axi_gmem_cout_RUSER;
input [1:0] m_axi_gmem_cout_RRESP;
input  m_axi_gmem_cout_BVALID;
output  m_axi_gmem_cout_BREADY;
input [1:0] m_axi_gmem_cout_BRESP;
input [1-1:0] m_axi_gmem_cout_BID;
input [1-1:0] m_axi_gmem_cout_BUSER;
input  ap_start;
output ap_done;
output ap_idle;
output ap_ready;
input  ap_continue;
input ap_clk;
input ap_rst_n;
(* keep_hierarchy = "yes" *)
kernel0_kernel0_gmem_cout_m_axi
#(
  .CONSERVATIVE(1),
  .USER_DW(512),
  .USER_AW(64),
  .USER_MAXREQS(5),
  .NUM_READ_OUTSTANDING(16),
  .NUM_WRITE_OUTSTANDING(16),
  .MAX_READ_BURST_LENGTH(16),
  .MAX_WRITE_BURST_LENGTH(16),
  .C_M_AXI_ID_WIDTH(C_M_AXI_GMEM_COUT_ID_WIDTH),
  .C_M_AXI_ADDR_WIDTH(C_M_AXI_GMEM_COUT_ADDR_WIDTH),
  .C_M_AXI_DATA_WIDTH(C_M_AXI_GMEM_COUT_DATA_WIDTH),
  .C_M_AXI_AWUSER_WIDTH(C_M_AXI_GMEM_COUT_AWUSER_WIDTH),
  .C_M_AXI_ARUSER_WIDTH(C_M_AXI_GMEM_COUT_ARUSER_WIDTH),
  .C_M_AXI_WUSER_WIDTH(C_M_AXI_GMEM_COUT_WUSER_WIDTH),
  .C_M_AXI_RUSER_WIDTH(C_M_AXI_GMEM_COUT_RUSER_WIDTH),
  .C_M_AXI_BUSER_WIDTH(C_M_AXI_GMEM_COUT_BUSER_WIDTH),
  .C_USER_VALUE(C_M_AXI_GMEM_COUT_USER_VALUE),
  .C_PROT_VALUE(C_M_AXI_GMEM_COUT_PROT_VALUE),
  .C_CACHE_VALUE(C_M_AXI_GMEM_COUT_CACHE_VALUE)
)
kernel0_gmem_cout_m_axi_U
(
  .AWVALID(m_axi_gmem_cout_AWVALID),
  .AWREADY(m_axi_gmem_cout_AWREADY),
  .AWADDR(m_axi_gmem_cout_AWADDR),
  .AWID(m_axi_gmem_cout_AWID),
  .AWLEN(m_axi_gmem_cout_AWLEN),
  .AWSIZE(m_axi_gmem_cout_AWSIZE),
  .AWBURST(m_axi_gmem_cout_AWBURST),
  .AWLOCK(m_axi_gmem_cout_AWLOCK),
  .AWCACHE(m_axi_gmem_cout_AWCACHE),
  .AWPROT(m_axi_gmem_cout_AWPROT),
  .AWQOS(m_axi_gmem_cout_AWQOS),
  .AWREGION(m_axi_gmem_cout_AWREGION),
  .AWUSER(m_axi_gmem_cout_AWUSER),
  .WVALID(m_axi_gmem_cout_WVALID),
  .WREADY(m_axi_gmem_cout_WREADY),
  .WDATA(m_axi_gmem_cout_WDATA),
  .WSTRB(m_axi_gmem_cout_WSTRB),
  .WLAST(m_axi_gmem_cout_WLAST),
  .WID(m_axi_gmem_cout_WID),
  .WUSER(m_axi_gmem_cout_WUSER),
  .ARVALID(m_axi_gmem_cout_ARVALID),
  .ARREADY(m_axi_gmem_cout_ARREADY),
  .ARADDR(m_axi_gmem_cout_ARADDR),
  .ARID(m_axi_gmem_cout_ARID),
  .ARLEN(m_axi_gmem_cout_ARLEN),
  .ARSIZE(m_axi_gmem_cout_ARSIZE),
  .ARBURST(m_axi_gmem_cout_ARBURST),
  .ARLOCK(m_axi_gmem_cout_ARLOCK),
  .ARCACHE(m_axi_gmem_cout_ARCACHE),
  .ARPROT(m_axi_gmem_cout_ARPROT),
  .ARQOS(m_axi_gmem_cout_ARQOS),
  .ARREGION(m_axi_gmem_cout_ARREGION),
  .ARUSER(m_axi_gmem_cout_ARUSER),
  .RVALID(m_axi_gmem_cout_RVALID),
  .RREADY(m_axi_gmem_cout_RREADY),
  .RDATA(m_axi_gmem_cout_RDATA),
  .RLAST(m_axi_gmem_cout_RLAST),
  .RID(m_axi_gmem_cout_RID),
  .RUSER(m_axi_gmem_cout_RUSER),
  .RRESP(m_axi_gmem_cout_RRESP),
  .BVALID(m_axi_gmem_cout_BVALID),
  .BREADY(m_axi_gmem_cout_BREADY),
  .BRESP(m_axi_gmem_cout_BRESP),
  .BID(m_axi_gmem_cout_BID),
  .BUSER(m_axi_gmem_cout_BUSER),
  .ACLK(ap_clk),
  .ARESET(ap_rst_pipe),
  .ACLK_EN(1'b1),
  .I_ARVALID(1'b0),
  .I_ARREADY(gmem_cout_ARREADY),
  .I_ARADDR(64'd0),
  .I_ARID(1'd0),
  .I_ARLEN(32'd0),
  .I_ARSIZE(3'd0),
  .I_ARLOCK(2'd0),
  .I_ARCACHE(4'd0),
  .I_ARQOS(4'd0),
  .I_ARPROT(3'd0),
  .I_ARUSER(1'd0),
  .I_ARBURST(2'd0),
  .I_ARREGION(4'd0),
  .I_RVALID(gmem_cout_RVALID),
  .I_RREADY(1'b0),
  .I_RDATA(gmem_cout_RDATA),
  .I_RID(gmem_cout_RID),
  .I_RUSER(gmem_cout_RUSER),
  .I_RRESP(gmem_cout_RRESP),
  .I_RLAST(gmem_cout_RLAST),
  .I_AWVALID(cout_drain_IO_L3_out_serialize_U0_m_axi_cout_V_AWVALID),
  .I_AWREADY(gmem_cout_AWREADY),
  .I_AWADDR(cout_drain_IO_L3_out_serialize_U0_m_axi_cout_V_AWADDR),
  .I_AWID(cout_drain_IO_L3_out_serialize_U0_m_axi_cout_V_AWID),
  .I_AWLEN(cout_drain_IO_L3_out_serialize_U0_m_axi_cout_V_AWLEN),
  .I_AWSIZE(cout_drain_IO_L3_out_serialize_U0_m_axi_cout_V_AWSIZE),
  .I_AWLOCK(cout_drain_IO_L3_out_serialize_U0_m_axi_cout_V_AWLOCK),
  .I_AWCACHE(cout_drain_IO_L3_out_serialize_U0_m_axi_cout_V_AWCACHE),
  .I_AWQOS(cout_drain_IO_L3_out_serialize_U0_m_axi_cout_V_AWQOS),
  .I_AWPROT(cout_drain_IO_L3_out_serialize_U0_m_axi_cout_V_AWPROT),
  .I_AWUSER(cout_drain_IO_L3_out_serialize_U0_m_axi_cout_V_AWUSER),
  .I_AWBURST(cout_drain_IO_L3_out_serialize_U0_m_axi_cout_V_AWBURST),
  .I_AWREGION(cout_drain_IO_L3_out_serialize_U0_m_axi_cout_V_AWREGION),
  .I_WVALID(cout_drain_IO_L3_out_serialize_U0_m_axi_cout_V_WVALID),
  .I_WREADY(gmem_cout_WREADY),
  .I_WDATA(cout_drain_IO_L3_out_serialize_U0_m_axi_cout_V_WDATA),
  .I_WID(cout_drain_IO_L3_out_serialize_U0_m_axi_cout_V_WID),
  .I_WUSER(cout_drain_IO_L3_out_serialize_U0_m_axi_cout_V_WUSER),
  .I_WLAST(cout_drain_IO_L3_out_serialize_U0_m_axi_cout_V_WLAST),
  .I_WSTRB(cout_drain_IO_L3_out_serialize_U0_m_axi_cout_V_WSTRB),
  .I_BVALID(gmem_cout_BVALID),
  .I_BREADY(cout_drain_IO_L3_out_serialize_U0_m_axi_cout_V_BREADY),
  .I_BRESP(gmem_cout_BRESP),
  .I_BID(gmem_cout_BID),
  .I_BUSER(gmem_cout_BUSER)
);

(* keep_hierarchy = "yes" *)
kernel0_PE_wrapper173
PE_wrapper173_U0
(
  .ap_clk(ap_clk),
  .ap_rst(ap_rst_pipe),
  .ap_start(ap_start_pipe),
  .ap_done(PE_wrapper173_U0_ap_done),
  .ap_continue(1'b1),
  .ap_idle(PE_wrapper173_U0_ap_idle),
  .ap_ready(PE_wrapper173_U0_ap_ready),
  .fifo_cin_in_V_V_dout(fifo_cin_PE_1_11_V_V_dout),
  .fifo_cin_in_V_V_empty_n(fifo_cin_PE_1_11_V_V_empty_n),
  .fifo_cin_in_V_V_read(PE_wrapper173_U0_fifo_cin_in_V_V_read),
  .fifo_cin_out_V_V_din(PE_wrapper173_U0_fifo_cin_out_V_V_din),
  .fifo_cin_out_V_V_full_n(fifo_cin_PE_2_11_V_V_full_n),
  .fifo_cin_out_V_V_write(PE_wrapper173_U0_fifo_cin_out_V_V_write),
  .fifo_cout_drain_out_V_din(PE_wrapper173_U0_fifo_cout_drain_out_V_din),
  .fifo_cout_drain_out_V_full_n(fifo_cout_drain_PE_1_11_V_full_n),
  .fifo_cout_drain_out_V_write(PE_wrapper173_U0_fifo_cout_drain_out_V_write),
  .fifo_w_in_V_V_dout(fifo_w_PE_1_11_V_V_dout),
  .fifo_w_in_V_V_empty_n(fifo_w_PE_1_11_V_V_empty_n),
  .fifo_w_in_V_V_read(PE_wrapper173_U0_fifo_w_in_V_V_read),
  .fifo_w_out_V_V_din(PE_wrapper173_U0_fifo_w_out_V_V_din),
  .fifo_w_out_V_V_full_n(fifo_w_PE_1_12_V_V_full_n),
  .fifo_w_out_V_V_write(PE_wrapper173_U0_fifo_w_out_V_V_write)
);

(* keep_hierarchy = "yes" *)
kernel0_PE_wrapper183
PE_wrapper183_U0
(
  .ap_clk(ap_clk),
  .ap_rst(ap_rst_pipe),
  .ap_start(ap_start_pipe),
  .ap_done(PE_wrapper183_U0_ap_done),
  .ap_continue(1'b1),
  .ap_idle(PE_wrapper183_U0_ap_idle),
  .ap_ready(PE_wrapper183_U0_ap_ready),
  .fifo_cin_in_V_V_dout(fifo_cin_PE_2_9_V_V_dout),
  .fifo_cin_in_V_V_empty_n(fifo_cin_PE_2_9_V_V_empty_n),
  .fifo_cin_in_V_V_read(PE_wrapper183_U0_fifo_cin_in_V_V_read),
  .fifo_cin_out_V_V_din(PE_wrapper183_U0_fifo_cin_out_V_V_din),
  .fifo_cin_out_V_V_full_n(fifo_cin_PE_3_9_V_V_full_n),
  .fifo_cin_out_V_V_write(PE_wrapper183_U0_fifo_cin_out_V_V_write),
  .fifo_cout_drain_out_V_din(PE_wrapper183_U0_fifo_cout_drain_out_V_din),
  .fifo_cout_drain_out_V_full_n(fifo_cout_drain_PE_2_9_V_full_n),
  .fifo_cout_drain_out_V_write(PE_wrapper183_U0_fifo_cout_drain_out_V_write),
  .fifo_w_in_V_V_dout(fifo_w_PE_2_9_V_V_dout),
  .fifo_w_in_V_V_empty_n(fifo_w_PE_2_9_V_V_empty_n),
  .fifo_w_in_V_V_read(PE_wrapper183_U0_fifo_w_in_V_V_read),
  .fifo_w_out_V_V_din(PE_wrapper183_U0_fifo_w_out_V_V_din),
  .fifo_w_out_V_V_full_n(fifo_w_PE_2_10_V_V_full_n),
  .fifo_w_out_V_V_write(PE_wrapper183_U0_fifo_w_out_V_V_write)
);

(* keep_hierarchy = "yes" *)
kernel0_PE_wrapper208
PE_wrapper208_U0
(
  .ap_clk(ap_clk),
  .ap_rst(ap_rst_pipe),
  .ap_start(ap_start_pipe),
  .ap_done(PE_wrapper208_U0_ap_done),
  .ap_continue(1'b1),
  .ap_idle(PE_wrapper208_U0_ap_idle),
  .ap_ready(PE_wrapper208_U0_ap_ready),
  .fifo_cin_in_V_V_dout(fifo_cin_PE_4_10_V_V_dout),
  .fifo_cin_in_V_V_empty_n(fifo_cin_PE_4_10_V_V_empty_n),
  .fifo_cin_in_V_V_read(PE_wrapper208_U0_fifo_cin_in_V_V_read),
  .fifo_cin_out_V_V_din(PE_wrapper208_U0_fifo_cin_out_V_V_din),
  .fifo_cin_out_V_V_full_n(fifo_cin_PE_5_10_V_V_full_n),
  .fifo_cin_out_V_V_write(PE_wrapper208_U0_fifo_cin_out_V_V_write),
  .fifo_cout_drain_out_V_din(PE_wrapper208_U0_fifo_cout_drain_out_V_din),
  .fifo_cout_drain_out_V_full_n(fifo_cout_drain_PE_4_10_V_full_n),
  .fifo_cout_drain_out_V_write(PE_wrapper208_U0_fifo_cout_drain_out_V_write),
  .fifo_w_in_V_V_dout(fifo_w_PE_4_10_V_V_dout),
  .fifo_w_in_V_V_empty_n(fifo_w_PE_4_10_V_V_empty_n),
  .fifo_w_in_V_V_read(PE_wrapper208_U0_fifo_w_in_V_V_read),
  .fifo_w_out_V_V_din(PE_wrapper208_U0_fifo_w_out_V_V_din),
  .fifo_w_out_V_V_full_n(fifo_w_PE_4_11_V_V_full_n),
  .fifo_w_out_V_V_write(PE_wrapper208_U0_fifo_w_out_V_V_write)
);

(* keep_hierarchy = "yes" *)
kernel0_PE_wrapper220
PE_wrapper220_U0
(
  .ap_clk(ap_clk),
  .ap_rst(ap_rst_pipe),
  .ap_start(ap_start_pipe),
  .ap_done(PE_wrapper220_U0_ap_done),
  .ap_continue(1'b1),
  .ap_idle(PE_wrapper220_U0_ap_idle),
  .ap_ready(PE_wrapper220_U0_ap_ready),
  .fifo_cin_in_V_V_dout(fifo_cin_PE_5_10_V_V_dout),
  .fifo_cin_in_V_V_empty_n(fifo_cin_PE_5_10_V_V_empty_n),
  .fifo_cin_in_V_V_read(PE_wrapper220_U0_fifo_cin_in_V_V_read),
  .fifo_cin_out_V_V_din(PE_wrapper220_U0_fifo_cin_out_V_V_din),
  .fifo_cin_out_V_V_full_n(fifo_cin_PE_6_10_V_V_full_n),
  .fifo_cin_out_V_V_write(PE_wrapper220_U0_fifo_cin_out_V_V_write),
  .fifo_cout_drain_out_V_din(PE_wrapper220_U0_fifo_cout_drain_out_V_din),
  .fifo_cout_drain_out_V_full_n(fifo_cout_drain_PE_5_10_V_full_n),
  .fifo_cout_drain_out_V_write(PE_wrapper220_U0_fifo_cout_drain_out_V_write),
  .fifo_w_in_V_V_dout(fifo_w_PE_5_10_V_V_dout),
  .fifo_w_in_V_V_empty_n(fifo_w_PE_5_10_V_V_empty_n),
  .fifo_w_in_V_V_read(PE_wrapper220_U0_fifo_w_in_V_V_read),
  .fifo_w_out_V_V_din(PE_wrapper220_U0_fifo_w_out_V_V_din),
  .fifo_w_out_V_V_full_n(fifo_w_PE_5_11_V_V_full_n),
  .fifo_w_out_V_V_write(PE_wrapper220_U0_fifo_w_out_V_V_write)
);

(* keep_hierarchy = "yes" *)
kernel0_PE_wrapper232
PE_wrapper232_U0
(
  .ap_clk(ap_clk),
  .ap_rst(ap_rst_pipe),
  .ap_start(ap_start_pipe),
  .ap_done(PE_wrapper232_U0_ap_done),
  .ap_continue(1'b1),
  .ap_idle(PE_wrapper232_U0_ap_idle),
  .ap_ready(PE_wrapper232_U0_ap_ready),
  .fifo_cin_in_V_V_dout(fifo_cin_PE_6_10_V_V_dout),
  .fifo_cin_in_V_V_empty_n(fifo_cin_PE_6_10_V_V_empty_n),
  .fifo_cin_in_V_V_read(PE_wrapper232_U0_fifo_cin_in_V_V_read),
  .fifo_cin_out_V_V_din(PE_wrapper232_U0_fifo_cin_out_V_V_din),
  .fifo_cin_out_V_V_full_n(fifo_cin_PE_7_10_V_V_full_n),
  .fifo_cin_out_V_V_write(PE_wrapper232_U0_fifo_cin_out_V_V_write),
  .fifo_cout_drain_out_V_din(PE_wrapper232_U0_fifo_cout_drain_out_V_din),
  .fifo_cout_drain_out_V_full_n(fifo_cout_drain_PE_6_10_V_full_n),
  .fifo_cout_drain_out_V_write(PE_wrapper232_U0_fifo_cout_drain_out_V_write),
  .fifo_w_in_V_V_dout(fifo_w_PE_6_10_V_V_dout),
  .fifo_w_in_V_V_empty_n(fifo_w_PE_6_10_V_V_empty_n),
  .fifo_w_in_V_V_read(PE_wrapper232_U0_fifo_w_in_V_V_read),
  .fifo_w_out_V_V_din(PE_wrapper232_U0_fifo_w_out_V_V_din),
  .fifo_w_out_V_V_full_n(fifo_w_PE_6_11_V_V_full_n),
  .fifo_w_out_V_V_write(PE_wrapper232_U0_fifo_w_out_V_V_write)
);

(* keep_hierarchy = "yes" *)
kernel0_PE_wrapper244
PE_wrapper244_U0
(
  .ap_clk(ap_clk),
  .ap_rst(ap_rst_pipe),
  .ap_start(ap_start_pipe),
  .ap_done(PE_wrapper244_U0_ap_done),
  .ap_continue(1'b1),
  .ap_idle(PE_wrapper244_U0_ap_idle),
  .ap_ready(PE_wrapper244_U0_ap_ready),
  .fifo_cin_in_V_V_dout(fifo_cin_PE_7_10_V_V_dout),
  .fifo_cin_in_V_V_empty_n(fifo_cin_PE_7_10_V_V_empty_n),
  .fifo_cin_in_V_V_read(PE_wrapper244_U0_fifo_cin_in_V_V_read),
  .fifo_cin_out_V_V_din(PE_wrapper244_U0_fifo_cin_out_V_V_din),
  .fifo_cin_out_V_V_full_n(fifo_cin_PE_8_10_V_V_full_n),
  .fifo_cin_out_V_V_write(PE_wrapper244_U0_fifo_cin_out_V_V_write),
  .fifo_cout_drain_out_V_din(PE_wrapper244_U0_fifo_cout_drain_out_V_din),
  .fifo_cout_drain_out_V_full_n(fifo_cout_drain_PE_7_10_V_full_n),
  .fifo_cout_drain_out_V_write(PE_wrapper244_U0_fifo_cout_drain_out_V_write),
  .fifo_w_in_V_V_dout(fifo_w_PE_7_10_V_V_dout),
  .fifo_w_in_V_V_empty_n(fifo_w_PE_7_10_V_V_empty_n),
  .fifo_w_in_V_V_read(PE_wrapper244_U0_fifo_w_in_V_V_read),
  .fifo_w_out_V_V_din(PE_wrapper244_U0_fifo_w_out_V_V_din),
  .fifo_w_out_V_V_full_n(fifo_w_PE_7_11_V_V_full_n),
  .fifo_w_out_V_V_write(PE_wrapper244_U0_fifo_w_out_V_V_write)
);

(* keep_hierarchy = "yes" *)
kernel0_PE_wrapper255
PE_wrapper255_U0
(
  .ap_clk(ap_clk),
  .ap_rst(ap_rst_pipe),
  .ap_start(ap_start_pipe),
  .ap_done(PE_wrapper255_U0_ap_done),
  .ap_continue(1'b1),
  .ap_idle(PE_wrapper255_U0_ap_idle),
  .ap_ready(PE_wrapper255_U0_ap_ready),
  .fifo_cin_in_V_V_dout(fifo_cin_PE_8_9_V_V_dout),
  .fifo_cin_in_V_V_empty_n(fifo_cin_PE_8_9_V_V_empty_n),
  .fifo_cin_in_V_V_read(PE_wrapper255_U0_fifo_cin_in_V_V_read),
  .fifo_cin_out_V_V_din(PE_wrapper255_U0_fifo_cin_out_V_V_din),
  .fifo_cin_out_V_V_full_n(fifo_cin_PE_9_9_V_V_full_n),
  .fifo_cin_out_V_V_write(PE_wrapper255_U0_fifo_cin_out_V_V_write),
  .fifo_cout_drain_out_V_din(PE_wrapper255_U0_fifo_cout_drain_out_V_din),
  .fifo_cout_drain_out_V_full_n(fifo_cout_drain_PE_8_9_V_full_n),
  .fifo_cout_drain_out_V_write(PE_wrapper255_U0_fifo_cout_drain_out_V_write),
  .fifo_w_in_V_V_dout(fifo_w_PE_8_9_V_V_dout),
  .fifo_w_in_V_V_empty_n(fifo_w_PE_8_9_V_V_empty_n),
  .fifo_w_in_V_V_read(PE_wrapper255_U0_fifo_w_in_V_V_read),
  .fifo_w_out_V_V_din(PE_wrapper255_U0_fifo_w_out_V_V_din),
  .fifo_w_out_V_V_full_n(fifo_w_PE_8_10_V_V_full_n),
  .fifo_w_out_V_V_write(PE_wrapper255_U0_fifo_w_out_V_V_write)
);

(* keep_hierarchy = "yes" *)
kernel0_w_PE_dummy_in357
w_PE_dummy_in357_U0
(
  .ap_clk(ap_clk),
  .ap_rst(ap_rst_pipe),
  .ap_start(ap_start_pipe),
  .ap_done(w_PE_dummy_in357_U0_ap_done),
  .ap_continue(1'b1),
  .ap_idle(w_PE_dummy_in357_U0_ap_idle),
  .ap_ready(w_PE_dummy_in357_U0_ap_ready),
  .fifo_w_in_V_V_dout(fifo_w_PE_5_12_V_V_dout),
  .fifo_w_in_V_V_empty_n(fifo_w_PE_5_12_V_V_empty_n),
  .fifo_w_in_V_V_read(w_PE_dummy_in357_U0_fifo_w_in_V_V_read)
);

(* keep_hierarchy = "yes" *)
kernel0_cout_drain_IO_L1_out_wrapper519
cout_drain_IO_L1_out_wrapper519_U0
(
  .ap_clk(ap_clk),
  .ap_rst(ap_rst_pipe),
  .ap_start(ap_start_pipe),
  .ap_done(cout_drain_IO_L1_out_wrapper519_U0_ap_done),
  .ap_continue(1'b1),
  .ap_idle(cout_drain_IO_L1_out_wrapper519_U0_ap_idle),
  .ap_ready(cout_drain_IO_L1_out_wrapper519_U0_ap_ready),
  .fifo_cout_drain_in_V_V_dout(fifo_cout_drain_cout_drain_IO_L1_out_9_8_V_V_dout),
  .fifo_cout_drain_in_V_V_empty_n(fifo_cout_drain_cout_drain_IO_L1_out_9_8_V_V_empty_n),
  .fifo_cout_drain_in_V_V_read(cout_drain_IO_L1_out_wrapper519_U0_fifo_cout_drain_in_V_V_read),
  .fifo_cout_drain_out_V_V_din(cout_drain_IO_L1_out_wrapper519_U0_fifo_cout_drain_out_V_V_din),
  .fifo_cout_drain_out_V_V_full_n(fifo_cout_drain_cout_drain_IO_L1_out_9_7_V_V_full_n),
  .fifo_cout_drain_out_V_V_write(cout_drain_IO_L1_out_wrapper519_U0_fifo_cout_drain_out_V_V_write),
  .fifo_cout_drain_local_in_V_dout(fifo_cout_drain_PE_7_9_V_dout),
  .fifo_cout_drain_local_in_V_empty_n(fifo_cout_drain_PE_7_9_V_empty_n),
  .fifo_cout_drain_local_in_V_read(cout_drain_IO_L1_out_wrapper519_U0_fifo_cout_drain_local_in_V_read)
);

(* keep_hierarchy = "yes" *)
kernel0_cout_drain_IO_L1_out_wrapper520
cout_drain_IO_L1_out_wrapper520_U0
(
  .ap_clk(ap_clk),
  .ap_rst(ap_rst_pipe),
  .ap_start(ap_start_pipe),
  .ap_done(cout_drain_IO_L1_out_wrapper520_U0_ap_done),
  .ap_continue(1'b1),
  .ap_idle(cout_drain_IO_L1_out_wrapper520_U0_ap_idle),
  .ap_ready(cout_drain_IO_L1_out_wrapper520_U0_ap_ready),
  .fifo_cout_drain_in_V_V_dout(fifo_cout_drain_cout_drain_IO_L1_out_9_7_V_V_dout),
  .fifo_cout_drain_in_V_V_empty_n(fifo_cout_drain_cout_drain_IO_L1_out_9_7_V_V_empty_n),
  .fifo_cout_drain_in_V_V_read(cout_drain_IO_L1_out_wrapper520_U0_fifo_cout_drain_in_V_V_read),
  .fifo_cout_drain_out_V_V_din(cout_drain_IO_L1_out_wrapper520_U0_fifo_cout_drain_out_V_V_din),
  .fifo_cout_drain_out_V_V_full_n(fifo_cout_drain_cout_drain_IO_L1_out_9_6_V_V_full_n),
  .fifo_cout_drain_out_V_V_write(cout_drain_IO_L1_out_wrapper520_U0_fifo_cout_drain_out_V_V_write),
  .fifo_cout_drain_local_in_V_dout(fifo_cout_drain_PE_6_9_V_dout),
  .fifo_cout_drain_local_in_V_empty_n(fifo_cout_drain_PE_6_9_V_empty_n),
  .fifo_cout_drain_local_in_V_read(cout_drain_IO_L1_out_wrapper520_U0_fifo_cout_drain_local_in_V_read)
);

(* keep_hierarchy = "yes" *)
kernel0_cout_drain_IO_L1_out_wrapper535
cout_drain_IO_L1_out_wrapper535_U0
(
  .ap_clk(ap_clk),
  .ap_rst(ap_rst_pipe),
  .ap_start(ap_start_pipe),
  .ap_done(cout_drain_IO_L1_out_wrapper535_U0_ap_done),
  .ap_continue(1'b1),
  .ap_idle(cout_drain_IO_L1_out_wrapper535_U0_ap_idle),
  .ap_ready(cout_drain_IO_L1_out_wrapper535_U0_ap_ready),
  .fifo_cout_drain_in_V_V_dout(fifo_cout_drain_cout_drain_IO_L1_out_10_8_V_V_dout),
  .fifo_cout_drain_in_V_V_empty_n(fifo_cout_drain_cout_drain_IO_L1_out_10_8_V_V_empty_n),
  .fifo_cout_drain_in_V_V_read(cout_drain_IO_L1_out_wrapper535_U0_fifo_cout_drain_in_V_V_read),
  .fifo_cout_drain_out_V_V_din(cout_drain_IO_L1_out_wrapper535_U0_fifo_cout_drain_out_V_V_din),
  .fifo_cout_drain_out_V_V_full_n(fifo_cout_drain_cout_drain_IO_L1_out_10_7_V_V_full_n),
  .fifo_cout_drain_out_V_V_write(cout_drain_IO_L1_out_wrapper535_U0_fifo_cout_drain_out_V_V_write),
  .fifo_cout_drain_local_in_V_dout(fifo_cout_drain_PE_7_10_V_dout),
  .fifo_cout_drain_local_in_V_empty_n(fifo_cout_drain_PE_7_10_V_empty_n),
  .fifo_cout_drain_local_in_V_read(cout_drain_IO_L1_out_wrapper535_U0_fifo_cout_drain_local_in_V_read)
);

(* keep_hierarchy = "yes" *)
kernel0_cout_drain_IO_L1_out_wrapper537
cout_drain_IO_L1_out_wrapper537_U0
(
  .ap_clk(ap_clk),
  .ap_rst(ap_rst_pipe),
  .ap_start(ap_start_pipe),
  .ap_done(cout_drain_IO_L1_out_wrapper537_U0_ap_done),
  .ap_continue(1'b1),
  .ap_idle(cout_drain_IO_L1_out_wrapper537_U0_ap_idle),
  .ap_ready(cout_drain_IO_L1_out_wrapper537_U0_ap_ready),
  .fifo_cout_drain_in_V_V_dout(fifo_cout_drain_cout_drain_IO_L1_out_10_6_V_V_dout),
  .fifo_cout_drain_in_V_V_empty_n(fifo_cout_drain_cout_drain_IO_L1_out_10_6_V_V_empty_n),
  .fifo_cout_drain_in_V_V_read(cout_drain_IO_L1_out_wrapper537_U0_fifo_cout_drain_in_V_V_read),
  .fifo_cout_drain_out_V_V_din(cout_drain_IO_L1_out_wrapper537_U0_fifo_cout_drain_out_V_V_din),
  .fifo_cout_drain_out_V_V_full_n(fifo_cout_drain_cout_drain_IO_L1_out_10_5_V_V_full_n),
  .fifo_cout_drain_out_V_V_write(cout_drain_IO_L1_out_wrapper537_U0_fifo_cout_drain_out_V_V_write),
  .fifo_cout_drain_local_in_V_dout(fifo_cout_drain_PE_5_10_V_dout),
  .fifo_cout_drain_local_in_V_empty_n(fifo_cout_drain_PE_5_10_V_empty_n),
  .fifo_cout_drain_local_in_V_read(cout_drain_IO_L1_out_wrapper537_U0_fifo_cout_drain_local_in_V_read)
);

(* keep_hierarchy = "yes" *)
kernel0_cout_drain_IO_L1_out_wrapper540
cout_drain_IO_L1_out_wrapper540_U0
(
  .ap_clk(ap_clk),
  .ap_rst(ap_rst_pipe),
  .ap_start(ap_start_pipe),
  .ap_done(cout_drain_IO_L1_out_wrapper540_U0_ap_done),
  .ap_continue(1'b1),
  .ap_idle(cout_drain_IO_L1_out_wrapper540_U0_ap_idle),
  .ap_ready(cout_drain_IO_L1_out_wrapper540_U0_ap_ready),
  .fifo_cout_drain_in_V_V_dout(fifo_cout_drain_cout_drain_IO_L1_out_10_3_V_V_dout),
  .fifo_cout_drain_in_V_V_empty_n(fifo_cout_drain_cout_drain_IO_L1_out_10_3_V_V_empty_n),
  .fifo_cout_drain_in_V_V_read(cout_drain_IO_L1_out_wrapper540_U0_fifo_cout_drain_in_V_V_read),
  .fifo_cout_drain_out_V_V_din(cout_drain_IO_L1_out_wrapper540_U0_fifo_cout_drain_out_V_V_din),
  .fifo_cout_drain_out_V_V_full_n(fifo_cout_drain_cout_drain_IO_L1_out_10_2_V_V_full_n),
  .fifo_cout_drain_out_V_V_write(cout_drain_IO_L1_out_wrapper540_U0_fifo_cout_drain_out_V_V_write),
  .fifo_cout_drain_local_in_V_dout(fifo_cout_drain_PE_2_10_V_dout),
  .fifo_cout_drain_local_in_V_empty_n(fifo_cout_drain_PE_2_10_V_empty_n),
  .fifo_cout_drain_local_in_V_read(cout_drain_IO_L1_out_wrapper540_U0_fifo_cout_drain_local_in_V_read)
);

(* keep_hierarchy = "yes" *)
kernel0_cout_drain_IO_L1_out_wrapper552
cout_drain_IO_L1_out_wrapper552_U0
(
  .ap_clk(ap_clk),
  .ap_rst(ap_rst_pipe),
  .ap_start(ap_start_pipe),
  .ap_done(cout_drain_IO_L1_out_wrapper552_U0_ap_done),
  .ap_continue(1'b1),
  .ap_idle(cout_drain_IO_L1_out_wrapper552_U0_ap_idle),
  .ap_ready(cout_drain_IO_L1_out_wrapper552_U0_ap_ready),
  .fifo_cout_drain_in_V_V_dout(fifo_cout_drain_cout_drain_IO_L1_out_11_6_V_V_dout),
  .fifo_cout_drain_in_V_V_empty_n(fifo_cout_drain_cout_drain_IO_L1_out_11_6_V_V_empty_n),
  .fifo_cout_drain_in_V_V_read(cout_drain_IO_L1_out_wrapper552_U0_fifo_cout_drain_in_V_V_read),
  .fifo_cout_drain_out_V_V_din(cout_drain_IO_L1_out_wrapper552_U0_fifo_cout_drain_out_V_V_din),
  .fifo_cout_drain_out_V_V_full_n(fifo_cout_drain_cout_drain_IO_L1_out_11_5_V_V_full_n),
  .fifo_cout_drain_out_V_V_write(cout_drain_IO_L1_out_wrapper552_U0_fifo_cout_drain_out_V_V_write),
  .fifo_cout_drain_local_in_V_dout(fifo_cout_drain_PE_5_11_V_dout),
  .fifo_cout_drain_local_in_V_empty_n(fifo_cout_drain_PE_5_11_V_empty_n),
  .fifo_cout_drain_local_in_V_read(cout_drain_IO_L1_out_wrapper552_U0_fifo_cout_drain_local_in_V_read)
);

(* keep_hierarchy = "yes" *)
kernel0_cout_drain_IO_L1_out_wrapper554
cout_drain_IO_L1_out_wrapper554_U0
(
  .ap_clk(ap_clk),
  .ap_rst(ap_rst_pipe),
  .ap_start(ap_start_pipe),
  .ap_done(cout_drain_IO_L1_out_wrapper554_U0_ap_done),
  .ap_continue(1'b1),
  .ap_idle(cout_drain_IO_L1_out_wrapper554_U0_ap_idle),
  .ap_ready(cout_drain_IO_L1_out_wrapper554_U0_ap_ready),
  .fifo_cout_drain_in_V_V_dout(fifo_cout_drain_cout_drain_IO_L1_out_11_4_V_V_dout),
  .fifo_cout_drain_in_V_V_empty_n(fifo_cout_drain_cout_drain_IO_L1_out_11_4_V_V_empty_n),
  .fifo_cout_drain_in_V_V_read(cout_drain_IO_L1_out_wrapper554_U0_fifo_cout_drain_in_V_V_read),
  .fifo_cout_drain_out_V_V_din(cout_drain_IO_L1_out_wrapper554_U0_fifo_cout_drain_out_V_V_din),
  .fifo_cout_drain_out_V_V_full_n(fifo_cout_drain_cout_drain_IO_L1_out_11_3_V_V_full_n),
  .fifo_cout_drain_out_V_V_write(cout_drain_IO_L1_out_wrapper554_U0_fifo_cout_drain_out_V_V_write),
  .fifo_cout_drain_local_in_V_dout(fifo_cout_drain_PE_3_11_V_dout),
  .fifo_cout_drain_local_in_V_empty_n(fifo_cout_drain_PE_3_11_V_empty_n),
  .fifo_cout_drain_local_in_V_read(cout_drain_IO_L1_out_wrapper554_U0_fifo_cout_drain_local_in_V_read)
);

(* keep_hierarchy = "yes" *)
kernel0_cout_drain_IO_L1_out_wrapper555
cout_drain_IO_L1_out_wrapper555_U0
(
  .ap_clk(ap_clk),
  .ap_rst(ap_rst_pipe),
  .ap_start(ap_start_pipe),
  .ap_done(cout_drain_IO_L1_out_wrapper555_U0_ap_done),
  .ap_continue(1'b1),
  .ap_idle(cout_drain_IO_L1_out_wrapper555_U0_ap_idle),
  .ap_ready(cout_drain_IO_L1_out_wrapper555_U0_ap_ready),
  .fifo_cout_drain_in_V_V_dout(fifo_cout_drain_cout_drain_IO_L1_out_11_3_V_V_dout),
  .fifo_cout_drain_in_V_V_empty_n(fifo_cout_drain_cout_drain_IO_L1_out_11_3_V_V_empty_n),
  .fifo_cout_drain_in_V_V_read(cout_drain_IO_L1_out_wrapper555_U0_fifo_cout_drain_in_V_V_read),
  .fifo_cout_drain_out_V_V_din(cout_drain_IO_L1_out_wrapper555_U0_fifo_cout_drain_out_V_V_din),
  .fifo_cout_drain_out_V_V_full_n(fifo_cout_drain_cout_drain_IO_L1_out_11_2_V_V_full_n),
  .fifo_cout_drain_out_V_V_write(cout_drain_IO_L1_out_wrapper555_U0_fifo_cout_drain_out_V_V_write),
  .fifo_cout_drain_local_in_V_dout(fifo_cout_drain_PE_2_11_V_dout),
  .fifo_cout_drain_local_in_V_empty_n(fifo_cout_drain_PE_2_11_V_empty_n),
  .fifo_cout_drain_local_in_V_read(cout_drain_IO_L1_out_wrapper555_U0_fifo_cout_drain_local_in_V_read)
);

(* keep_hierarchy = "yes" *)
kernel0_cout_drain_IO_L3_out_serialize
cout_drain_IO_L3_out_serialize_U0
(
  .ap_clk(ap_clk),
  .ap_rst(ap_rst_pipe),
  .ap_start(ap_start_pipe),
  .ap_done(cout_drain_IO_L3_out_serialize_U0_ap_done),
  .ap_continue(1'b1),
  .ap_idle(cout_drain_IO_L3_out_serialize_U0_ap_idle),
  .ap_ready(cout_drain_IO_L3_out_serialize_U0_ap_ready),
  .m_axi_cout_V_AWVALID(cout_drain_IO_L3_out_serialize_U0_m_axi_cout_V_AWVALID),
  .m_axi_cout_V_AWREADY(gmem_cout_AWREADY),
  .m_axi_cout_V_AWADDR(cout_drain_IO_L3_out_serialize_U0_m_axi_cout_V_AWADDR),
  .m_axi_cout_V_AWID(cout_drain_IO_L3_out_serialize_U0_m_axi_cout_V_AWID),
  .m_axi_cout_V_AWLEN(cout_drain_IO_L3_out_serialize_U0_m_axi_cout_V_AWLEN),
  .m_axi_cout_V_AWSIZE(cout_drain_IO_L3_out_serialize_U0_m_axi_cout_V_AWSIZE),
  .m_axi_cout_V_AWBURST(cout_drain_IO_L3_out_serialize_U0_m_axi_cout_V_AWBURST),
  .m_axi_cout_V_AWLOCK(cout_drain_IO_L3_out_serialize_U0_m_axi_cout_V_AWLOCK),
  .m_axi_cout_V_AWCACHE(cout_drain_IO_L3_out_serialize_U0_m_axi_cout_V_AWCACHE),
  .m_axi_cout_V_AWPROT(cout_drain_IO_L3_out_serialize_U0_m_axi_cout_V_AWPROT),
  .m_axi_cout_V_AWQOS(cout_drain_IO_L3_out_serialize_U0_m_axi_cout_V_AWQOS),
  .m_axi_cout_V_AWREGION(cout_drain_IO_L3_out_serialize_U0_m_axi_cout_V_AWREGION),
  .m_axi_cout_V_AWUSER(cout_drain_IO_L3_out_serialize_U0_m_axi_cout_V_AWUSER),
  .m_axi_cout_V_WVALID(cout_drain_IO_L3_out_serialize_U0_m_axi_cout_V_WVALID),
  .m_axi_cout_V_WREADY(gmem_cout_WREADY),
  .m_axi_cout_V_WDATA(cout_drain_IO_L3_out_serialize_U0_m_axi_cout_V_WDATA),
  .m_axi_cout_V_WSTRB(cout_drain_IO_L3_out_serialize_U0_m_axi_cout_V_WSTRB),
  .m_axi_cout_V_WLAST(cout_drain_IO_L3_out_serialize_U0_m_axi_cout_V_WLAST),
  .m_axi_cout_V_WID(cout_drain_IO_L3_out_serialize_U0_m_axi_cout_V_WID),
  .m_axi_cout_V_WUSER(cout_drain_IO_L3_out_serialize_U0_m_axi_cout_V_WUSER),
  .m_axi_cout_V_ARVALID(cout_drain_IO_L3_out_serialize_U0_m_axi_cout_V_ARVALID),
  .m_axi_cout_V_ARREADY(1'b0),
  .m_axi_cout_V_ARADDR(cout_drain_IO_L3_out_serialize_U0_m_axi_cout_V_ARADDR),
  .m_axi_cout_V_ARID(cout_drain_IO_L3_out_serialize_U0_m_axi_cout_V_ARID),
  .m_axi_cout_V_ARLEN(cout_drain_IO_L3_out_serialize_U0_m_axi_cout_V_ARLEN),
  .m_axi_cout_V_ARSIZE(cout_drain_IO_L3_out_serialize_U0_m_axi_cout_V_ARSIZE),
  .m_axi_cout_V_ARBURST(cout_drain_IO_L3_out_serialize_U0_m_axi_cout_V_ARBURST),
  .m_axi_cout_V_ARLOCK(cout_drain_IO_L3_out_serialize_U0_m_axi_cout_V_ARLOCK),
  .m_axi_cout_V_ARCACHE(cout_drain_IO_L3_out_serialize_U0_m_axi_cout_V_ARCACHE),
  .m_axi_cout_V_ARPROT(cout_drain_IO_L3_out_serialize_U0_m_axi_cout_V_ARPROT),
  .m_axi_cout_V_ARQOS(cout_drain_IO_L3_out_serialize_U0_m_axi_cout_V_ARQOS),
  .m_axi_cout_V_ARREGION(cout_drain_IO_L3_out_serialize_U0_m_axi_cout_V_ARREGION),
  .m_axi_cout_V_ARUSER(cout_drain_IO_L3_out_serialize_U0_m_axi_cout_V_ARUSER),
  .m_axi_cout_V_RVALID(1'b0),
  .m_axi_cout_V_RREADY(cout_drain_IO_L3_out_serialize_U0_m_axi_cout_V_RREADY),
  .m_axi_cout_V_RDATA(512'd0),
  .m_axi_cout_V_RLAST(1'b0),
  .m_axi_cout_V_RID(1'd0),
  .m_axi_cout_V_RUSER(1'd0),
  .m_axi_cout_V_RRESP(2'd0),
  .m_axi_cout_V_BVALID(gmem_cout_BVALID),
  .m_axi_cout_V_BREADY(cout_drain_IO_L3_out_serialize_U0_m_axi_cout_V_BREADY),
  .m_axi_cout_V_BRESP(gmem_cout_BRESP),
  .m_axi_cout_V_BID(gmem_cout_BID),
  .m_axi_cout_V_BUSER(gmem_cout_BUSER),
  .cout_V_offset_dout(cout_V_c_dout),
  .cout_V_offset_empty_n(cout_V_c_empty_n),
  .cout_V_offset_read(cout_drain_IO_L3_out_serialize_U0_cout_V_offset_read),
  .fifo_cout_drain_local_in_V_V_dout(fifo_cout_drain_cout_drain_IO_L3_out_serialize_V_V_dout),
  .fifo_cout_drain_local_in_V_V_empty_n(fifo_cout_drain_cout_drain_IO_L3_out_serialize_V_V_empty_n),
  .fifo_cout_drain_local_in_V_V_read(cout_drain_IO_L3_out_serialize_U0_fifo_cout_drain_local_in_V_V_read)
);

(* keep_hierarchy = "yes" *)
fifo_almost_full
#(
  .DATA_WIDTH(256),
  .DEPTH(11),
  .ADDR_WIDTH(9),
  .GRACE_PERIOD(1)
)
fifo_cin_PE_7_10_V_V_U
(
  .clk(ap_clk),
  .reset(ap_rst_n_inv),
  .if_read_ce(1'b1),
  .if_write_ce(1'b1),
  .if_din(PE_wrapper232_U0_fifo_cin_out_V_V_din),
  .if_full_n(fifo_cin_PE_7_10_V_V_full_n),
  .if_write(PE_wrapper232_U0_fifo_cin_out_V_V_write),
  .if_dout(fifo_cin_PE_7_10_V_V_dout),
  .if_empty_n(fifo_cin_PE_7_10_V_V_empty_n),
  .if_read(PE_wrapper244_U0_fifo_cin_in_V_V_read)
);

(* keep_hierarchy = "yes" *)
fifo_almost_full
#(
  .DATA_WIDTH(32),
  .DEPTH(33),
  .ADDR_WIDTH(6),
  .GRACE_PERIOD(1)
)
fifo_cout_drain_PE_7_10_V_U
(
  .clk(ap_clk),
  .reset(ap_rst_n_inv),
  .if_read_ce(1'b1),
  .if_write_ce(1'b1),
  .if_din(PE_wrapper244_U0_fifo_cout_drain_out_V_din),
  .if_full_n(fifo_cout_drain_PE_7_10_V_full_n),
  .if_write(PE_wrapper244_U0_fifo_cout_drain_out_V_write),
  .if_dout(fifo_cout_drain_PE_7_10_V_dout),
  .if_empty_n(fifo_cout_drain_PE_7_10_V_empty_n),
  .if_read(cout_drain_IO_L1_out_wrapper535_U0_fifo_cout_drain_local_in_V_read)
);

(* keep_hierarchy = "yes" *)
fifo_almost_full
#(
  .DATA_WIDTH(64),
  .DEPTH(3),
  .ADDR_WIDTH(7),
  .GRACE_PERIOD(1)
)
fifo_cout_drain_cout_drain_IO_L1_out_11_3_V_V_U
(
  .clk(ap_clk),
  .reset(ap_rst_n_inv),
  .if_read_ce(1'b1),
  .if_write_ce(1'b1),
  .if_din(cout_drain_IO_L1_out_wrapper554_U0_fifo_cout_drain_out_V_V_din),
  .if_full_n(fifo_cout_drain_cout_drain_IO_L1_out_11_3_V_V_full_n),
  .if_write(cout_drain_IO_L1_out_wrapper554_U0_fifo_cout_drain_out_V_V_write),
  .if_dout(fifo_cout_drain_cout_drain_IO_L1_out_11_3_V_V_dout),
  .if_empty_n(fifo_cout_drain_cout_drain_IO_L1_out_11_3_V_V_empty_n),
  .if_read(cout_drain_IO_L1_out_wrapper555_U0_fifo_cout_drain_in_V_V_read)
);

(* keep_hierarchy = "yes" *)
fifo_almost_full
#(
  .DATA_WIDTH(32),
  .DEPTH(49),
  .ADDR_WIDTH(6),
  .GRACE_PERIOD(1)
)
fifo_cout_drain_PE_5_10_V_U
(
  .clk(ap_clk),
  .reset(ap_rst_n_inv),
  .if_read_ce(1'b1),
  .if_write_ce(1'b1),
  .if_din(PE_wrapper220_U0_fifo_cout_drain_out_V_din),
  .if_full_n(fifo_cout_drain_PE_5_10_V_full_n),
  .if_write(PE_wrapper220_U0_fifo_cout_drain_out_V_write),
  .if_dout(fifo_cout_drain_PE_5_10_V_dout),
  .if_empty_n(fifo_cout_drain_PE_5_10_V_empty_n),
  .if_read(cout_drain_IO_L1_out_wrapper537_U0_fifo_cout_drain_local_in_V_read)
);

(* keep_hierarchy = "yes" *)
fifo_almost_full
#(
  .DATA_WIDTH(256),
  .DEPTH(3),
  .ADDR_WIDTH(9),
  .GRACE_PERIOD(1)
)
fifo_cin_PE_5_10_V_V_U
(
  .clk(ap_clk),
  .reset(ap_rst_n_inv),
  .if_read_ce(1'b1),
  .if_write_ce(1'b1),
  .if_din(PE_wrapper208_U0_fifo_cin_out_V_V_din),
  .if_full_n(fifo_cin_PE_5_10_V_V_full_n),
  .if_write(PE_wrapper208_U0_fifo_cin_out_V_V_write),
  .if_dout(fifo_cin_PE_5_10_V_V_dout),
  .if_empty_n(fifo_cin_PE_5_10_V_V_empty_n),
  .if_read(PE_wrapper220_U0_fifo_cin_in_V_V_read)
);

(* keep_hierarchy = "yes" *)
fifo_almost_full
#(
  .DATA_WIDTH(64),
  .DEPTH(3),
  .ADDR_WIDTH(7),
  .GRACE_PERIOD(1)
)
fifo_cout_drain_cout_drain_IO_L1_out_9_7_V_V_U
(
  .clk(ap_clk),
  .reset(ap_rst_n_inv),
  .if_read_ce(1'b1),
  .if_write_ce(1'b1),
  .if_din(cout_drain_IO_L1_out_wrapper519_U0_fifo_cout_drain_out_V_V_din),
  .if_full_n(fifo_cout_drain_cout_drain_IO_L1_out_9_7_V_V_full_n),
  .if_write(cout_drain_IO_L1_out_wrapper519_U0_fifo_cout_drain_out_V_V_write),
  .if_dout(fifo_cout_drain_cout_drain_IO_L1_out_9_7_V_V_dout),
  .if_empty_n(fifo_cout_drain_cout_drain_IO_L1_out_9_7_V_V_empty_n),
  .if_read(cout_drain_IO_L1_out_wrapper520_U0_fifo_cout_drain_in_V_V_read)
);

(* keep_hierarchy = "yes" *)
fifo_almost_full
#(
  .DATA_WIDTH(256),
  .DEPTH(5),
  .ADDR_WIDTH(9),
  .GRACE_PERIOD(1)
)
fifo_cin_PE_6_10_V_V_U
(
  .clk(ap_clk),
  .reset(ap_rst_n_inv),
  .if_read_ce(1'b1),
  .if_write_ce(1'b1),
  .if_din(PE_wrapper220_U0_fifo_cin_out_V_V_din),
  .if_full_n(fifo_cin_PE_6_10_V_V_full_n),
  .if_write(PE_wrapper220_U0_fifo_cin_out_V_V_write),
  .if_dout(fifo_cin_PE_6_10_V_V_dout),
  .if_empty_n(fifo_cin_PE_6_10_V_V_empty_n),
  .if_read(PE_wrapper232_U0_fifo_cin_in_V_V_read)
);

(* keep_hierarchy = "yes" *)
fifo_almost_full
#(
  .DATA_WIDTH(256),
  .DEPTH(4),
  .ADDR_WIDTH(9),
  .GRACE_PERIOD(3)
)
fifo_w_PE_5_10_V_V_U
(
  .clk(ap_clk),
  .reset(ap_rst_n_inv),
  .if_read_ce(1'b1),
  .if_write_ce(1'b1),
  .if_din(PE_wrapper219_U0_fifo_w_out_V_V_din),
  .if_full_n(fifo_w_PE_5_10_V_V_full_n),
  .if_write(PE_wrapper219_U0_fifo_w_out_V_V_write),
  .if_dout(fifo_w_PE_5_10_V_V_dout),
  .if_empty_n(fifo_w_PE_5_10_V_V_empty_n),
  .if_read(PE_wrapper220_U0_fifo_w_in_V_V_read)
);

(* keep_hierarchy = "yes" *)
fifo_almost_full
#(
  .DATA_WIDTH(256),
  .DEPTH(4),
  .ADDR_WIDTH(9),
  .GRACE_PERIOD(3)
)
fifo_cin_PE_2_9_V_V_U
(
  .clk(ap_clk),
  .reset(ap_rst_n_inv),
  .if_read_ce(1'b1),
  .if_write_ce(1'b1),
  .if_din(PE_wrapper171_U0_fifo_cin_out_V_V_din),
  .if_full_n(fifo_cin_PE_2_9_V_V_full_n),
  .if_write(PE_wrapper171_U0_fifo_cin_out_V_V_write),
  .if_dout(fifo_cin_PE_2_9_V_V_dout),
  .if_empty_n(fifo_cin_PE_2_9_V_V_empty_n),
  .if_read(PE_wrapper183_U0_fifo_cin_in_V_V_read)
);

(* keep_hierarchy = "yes" *)
fifo_almost_full
#(
  .DATA_WIDTH(256),
  .DEPTH(4),
  .ADDR_WIDTH(9),
  .GRACE_PERIOD(3)
)
fifo_w_PE_1_11_V_V_U
(
  .clk(ap_clk),
  .reset(ap_rst_n_inv),
  .if_read_ce(1'b1),
  .if_write_ce(1'b1),
  .if_din(PE_wrapper172_U0_fifo_w_out_V_V_din),
  .if_full_n(fifo_w_PE_1_11_V_V_full_n),
  .if_write(PE_wrapper172_U0_fifo_w_out_V_V_write),
  .if_dout(fifo_w_PE_1_11_V_V_dout),
  .if_empty_n(fifo_w_PE_1_11_V_V_empty_n),
  .if_read(PE_wrapper173_U0_fifo_w_in_V_V_read)
);

(* keep_hierarchy = "yes" *)
fifo_almost_full
#(
  .DATA_WIDTH(64),
  .DEPTH(5),
  .ADDR_WIDTH(7),
  .GRACE_PERIOD(5)
)
fifo_cout_drain_cout_drain_IO_L1_out_11_6_V_V_U
(
  .clk(ap_clk),
  .reset(ap_rst_n_inv),
  .if_read_ce(1'b1),
  .if_write_ce(1'b1),
  .if_din(cout_drain_IO_L1_out_wrapper551_U0_fifo_cout_drain_out_V_V_din),
  .if_full_n(fifo_cout_drain_cout_drain_IO_L1_out_11_6_V_V_full_n),
  .if_write(cout_drain_IO_L1_out_wrapper551_U0_fifo_cout_drain_out_V_V_write),
  .if_dout(fifo_cout_drain_cout_drain_IO_L1_out_11_6_V_V_dout),
  .if_empty_n(fifo_cout_drain_cout_drain_IO_L1_out_11_6_V_V_empty_n),
  .if_read(cout_drain_IO_L1_out_wrapper552_U0_fifo_cout_drain_in_V_V_read)
);

(* keep_hierarchy = "yes" *)
fifo_almost_full
#(
  .DATA_WIDTH(256),
  .DEPTH(4),
  .ADDR_WIDTH(9),
  .GRACE_PERIOD(3)
)
fifo_cin_PE_4_10_V_V_U
(
  .clk(ap_clk),
  .reset(ap_rst_n_inv),
  .if_read_ce(1'b1),
  .if_write_ce(1'b1),
  .if_din(PE_wrapper196_U0_fifo_cin_out_V_V_din),
  .if_full_n(fifo_cin_PE_4_10_V_V_full_n),
  .if_write(PE_wrapper196_U0_fifo_cin_out_V_V_write),
  .if_dout(fifo_cin_PE_4_10_V_V_dout),
  .if_empty_n(fifo_cin_PE_4_10_V_V_empty_n),
  .if_read(PE_wrapper208_U0_fifo_cin_in_V_V_read)
);

(* keep_hierarchy = "yes" *)
fifo_almost_full
#(
  .DATA_WIDTH(64),
  .DEPTH(4),
  .ADDR_WIDTH(7),
  .GRACE_PERIOD(3)
)
fifo_cout_drain_cout_drain_IO_L1_out_10_3_V_V_U
(
  .clk(ap_clk),
  .reset(ap_rst_n_inv),
  .if_read_ce(1'b1),
  .if_write_ce(1'b1),
  .if_din(cout_drain_IO_L1_out_wrapper539_U0_fifo_cout_drain_out_V_V_din),
  .if_full_n(fifo_cout_drain_cout_drain_IO_L1_out_10_3_V_V_full_n),
  .if_write(cout_drain_IO_L1_out_wrapper539_U0_fifo_cout_drain_out_V_V_write),
  .if_dout(fifo_cout_drain_cout_drain_IO_L1_out_10_3_V_V_dout),
  .if_empty_n(fifo_cout_drain_cout_drain_IO_L1_out_10_3_V_V_empty_n),
  .if_read(cout_drain_IO_L1_out_wrapper540_U0_fifo_cout_drain_in_V_V_read)
);

(* keep_hierarchy = "yes" *)
fifo_almost_full
#(
  .DATA_WIDTH(256),
  .DEPTH(4),
  .ADDR_WIDTH(9),
  .GRACE_PERIOD(3)
)
fifo_w_PE_6_10_V_V_U
(
  .clk(ap_clk),
  .reset(ap_rst_n_inv),
  .if_read_ce(1'b1),
  .if_write_ce(1'b1),
  .if_din(PE_wrapper231_U0_fifo_w_out_V_V_din),
  .if_full_n(fifo_w_PE_6_10_V_V_full_n),
  .if_write(PE_wrapper231_U0_fifo_w_out_V_V_write),
  .if_dout(fifo_w_PE_6_10_V_V_dout),
  .if_empty_n(fifo_w_PE_6_10_V_V_empty_n),
  .if_read(PE_wrapper232_U0_fifo_w_in_V_V_read)
);

(* keep_hierarchy = "yes" *)
fifo_almost_full
#(
  .DATA_WIDTH(32),
  .DEPTH(40),
  .ADDR_WIDTH(6),
  .GRACE_PERIOD(3)
)
fifo_cout_drain_PE_6_9_V_U
(
  .clk(ap_clk),
  .reset(ap_rst_n_inv),
  .if_read_ce(1'b1),
  .if_write_ce(1'b1),
  .if_din(PE_wrapper231_U0_fifo_cout_drain_out_V_din),
  .if_full_n(fifo_cout_drain_PE_6_9_V_full_n),
  .if_write(PE_wrapper231_U0_fifo_cout_drain_out_V_write),
  .if_dout(fifo_cout_drain_PE_6_9_V_dout),
  .if_empty_n(fifo_cout_drain_PE_6_9_V_empty_n),
  .if_read(cout_drain_IO_L1_out_wrapper520_U0_fifo_cout_drain_local_in_V_read)
);

(* keep_hierarchy = "yes" *)
fifo_almost_full
#(
  .DATA_WIDTH(256),
  .DEPTH(4),
  .ADDR_WIDTH(9),
  .GRACE_PERIOD(3)
)
fifo_w_PE_4_10_V_V_U
(
  .clk(ap_clk),
  .reset(ap_rst_n_inv),
  .if_read_ce(1'b1),
  .if_write_ce(1'b1),
  .if_din(PE_wrapper207_U0_fifo_w_out_V_V_din),
  .if_full_n(fifo_w_PE_4_10_V_V_full_n),
  .if_write(PE_wrapper207_U0_fifo_w_out_V_V_write),
  .if_dout(fifo_w_PE_4_10_V_V_dout),
  .if_empty_n(fifo_w_PE_4_10_V_V_empty_n),
  .if_read(PE_wrapper208_U0_fifo_w_in_V_V_read)
);

(* keep_hierarchy = "yes" *)
fifo_almost_full
#(
  .DATA_WIDTH(32),
  .DEPTH(46),
  .ADDR_WIDTH(6),
  .GRACE_PERIOD(3)
)
fifo_cout_drain_PE_5_11_V_U
(
  .clk(ap_clk),
  .reset(ap_rst_n_inv),
  .if_read_ce(1'b1),
  .if_write_ce(1'b1),
  .if_din(PE_wrapper221_U0_fifo_cout_drain_out_V_din),
  .if_full_n(fifo_cout_drain_PE_5_11_V_full_n),
  .if_write(PE_wrapper221_U0_fifo_cout_drain_out_V_write),
  .if_dout(fifo_cout_drain_PE_5_11_V_dout),
  .if_empty_n(fifo_cout_drain_PE_5_11_V_empty_n),
  .if_read(cout_drain_IO_L1_out_wrapper552_U0_fifo_cout_drain_local_in_V_read)
);

(* keep_hierarchy = "yes" *)
fifo_almost_full
#(
  .DATA_WIDTH(256),
  .DEPTH(5),
  .ADDR_WIDTH(9),
  .GRACE_PERIOD(5)
)
fifo_cin_PE_1_11_V_V_U
(
  .clk(ap_clk),
  .reset(ap_rst_n_inv),
  .if_read_ce(1'b1),
  .if_write_ce(1'b1),
  .if_din(PE_wrapper161_U0_fifo_cin_out_V_V_din),
  .if_full_n(fifo_cin_PE_1_11_V_V_full_n),
  .if_write(PE_wrapper161_U0_fifo_cin_out_V_V_write),
  .if_dout(fifo_cin_PE_1_11_V_V_dout),
  .if_empty_n(fifo_cin_PE_1_11_V_V_empty_n),
  .if_read(PE_wrapper173_U0_fifo_cin_in_V_V_read)
);

(* keep_hierarchy = "yes" *)
fifo_almost_full
#(
  .DATA_WIDTH(64),
  .DEPTH(189),
  .ADDR_WIDTH(7),
  .GRACE_PERIOD(13)
)
cout_V_c_U
(
  .clk(ap_clk),
  .reset(ap_rst_n_inv),
  .if_read_ce(1'b1),
  .if_write_ce(1'b1),
  .if_din(kernel0_entry12_U0_cout_V_out_din),
  .if_full_n(cout_V_c_full_n),
  .if_write(kernel0_entry12_U0_cout_V_out_write),
  .if_dout(cout_V_c_dout),
  .if_empty_n(cout_V_c_empty_n),
  .if_read(cout_drain_IO_L3_out_serialize_U0_cout_V_offset_read)
);

(* keep_hierarchy = "yes" *)
fifo_almost_full
#(
  .DATA_WIDTH(256),
  .DEPTH(7),
  .ADDR_WIDTH(9),
  .GRACE_PERIOD(9)
)
fifo_w_PE_7_10_V_V_U
(
  .clk(ap_clk),
  .reset(ap_rst_n_inv),
  .if_read_ce(1'b1),
  .if_write_ce(1'b1),
  .if_din(PE_wrapper243_U0_fifo_w_out_V_V_din),
  .if_full_n(fifo_w_PE_7_10_V_V_full_n),
  .if_write(PE_wrapper243_U0_fifo_w_out_V_V_write),
  .if_dout(fifo_w_PE_7_10_V_V_dout),
  .if_empty_n(fifo_w_PE_7_10_V_V_empty_n),
  .if_read(PE_wrapper244_U0_fifo_w_in_V_V_read)
);

(* keep_hierarchy = "yes" *)
fifo_almost_full
#(
  .DATA_WIDTH(32),
  .DEPTH(33),
  .ADDR_WIDTH(6),
  .GRACE_PERIOD(9)
)
fifo_cout_drain_PE_7_9_V_U
(
  .clk(ap_clk),
  .reset(ap_rst_n_inv),
  .if_read_ce(1'b1),
  .if_write_ce(1'b1),
  .if_din(PE_wrapper243_U0_fifo_cout_drain_out_V_din),
  .if_full_n(fifo_cout_drain_PE_7_9_V_full_n),
  .if_write(PE_wrapper243_U0_fifo_cout_drain_out_V_write),
  .if_dout(fifo_cout_drain_PE_7_9_V_dout),
  .if_empty_n(fifo_cout_drain_PE_7_9_V_empty_n),
  .if_read(cout_drain_IO_L1_out_wrapper519_U0_fifo_cout_drain_local_in_V_read)
);

(* keep_hierarchy = "yes" *)
fifo_almost_full
#(
  .DATA_WIDTH(32),
  .DEPTH(58),
  .ADDR_WIDTH(6),
  .GRACE_PERIOD(3)
)
fifo_cout_drain_PE_2_10_V_U
(
  .clk(ap_clk),
  .reset(ap_rst_n_inv),
  .if_read_ce(1'b1),
  .if_write_ce(1'b1),
  .if_din(PE_wrapper184_U0_fifo_cout_drain_out_V_din),
  .if_full_n(fifo_cout_drain_PE_2_10_V_full_n),
  .if_write(PE_wrapper184_U0_fifo_cout_drain_out_V_write),
  .if_dout(fifo_cout_drain_PE_2_10_V_dout),
  .if_empty_n(fifo_cout_drain_PE_2_10_V_empty_n),
  .if_read(cout_drain_IO_L1_out_wrapper540_U0_fifo_cout_drain_local_in_V_read)
);

(* keep_hierarchy = "yes" *)
fifo_almost_full
#(
  .DATA_WIDTH(256),
  .DEPTH(7),
  .ADDR_WIDTH(9),
  .GRACE_PERIOD(9)
)
fifo_cin_PE_8_9_V_V_U
(
  .clk(ap_clk),
  .reset(ap_rst_n_inv),
  .if_read_ce(1'b1),
  .if_write_ce(1'b1),
  .if_din(PE_wrapper243_U0_fifo_cin_out_V_V_din),
  .if_full_n(fifo_cin_PE_8_9_V_V_full_n),
  .if_write(PE_wrapper243_U0_fifo_cin_out_V_V_write),
  .if_dout(fifo_cin_PE_8_9_V_V_dout),
  .if_empty_n(fifo_cin_PE_8_9_V_V_empty_n),
  .if_read(PE_wrapper255_U0_fifo_cin_in_V_V_read)
);

(* keep_hierarchy = "yes" *)
fifo_almost_full
#(
  .DATA_WIDTH(32),
  .DEPTH(55),
  .ADDR_WIDTH(6),
  .GRACE_PERIOD(5)
)
fifo_cout_drain_PE_2_11_V_U
(
  .clk(ap_clk),
  .reset(ap_rst_n_inv),
  .if_read_ce(1'b1),
  .if_write_ce(1'b1),
  .if_din(PE_wrapper185_U0_fifo_cout_drain_out_V_din),
  .if_full_n(fifo_cout_drain_PE_2_11_V_full_n),
  .if_write(PE_wrapper185_U0_fifo_cout_drain_out_V_write),
  .if_dout(fifo_cout_drain_PE_2_11_V_dout),
  .if_empty_n(fifo_cout_drain_PE_2_11_V_empty_n),
  .if_read(cout_drain_IO_L1_out_wrapper555_U0_fifo_cout_drain_local_in_V_read)
);

(* keep_hierarchy = "yes" *)
fifo_almost_full
#(
  .DATA_WIDTH(64),
  .DEPTH(5),
  .ADDR_WIDTH(7),
  .GRACE_PERIOD(5)
)
fifo_cout_drain_cout_drain_IO_L1_out_9_8_V_V_U
(
  .clk(ap_clk),
  .reset(ap_rst_n_inv),
  .if_read_ce(1'b1),
  .if_write_ce(1'b1),
  .if_din(cout_drain_IO_L1_out_wrapper518_U0_fifo_cout_drain_out_V_V_din),
  .if_full_n(fifo_cout_drain_cout_drain_IO_L1_out_9_8_V_V_full_n),
  .if_write(cout_drain_IO_L1_out_wrapper518_U0_fifo_cout_drain_out_V_V_write),
  .if_dout(fifo_cout_drain_cout_drain_IO_L1_out_9_8_V_V_dout),
  .if_empty_n(fifo_cout_drain_cout_drain_IO_L1_out_9_8_V_V_empty_n),
  .if_read(cout_drain_IO_L1_out_wrapper519_U0_fifo_cout_drain_in_V_V_read)
);

(* keep_hierarchy = "yes" *)
fifo_almost_full
#(
  .DATA_WIDTH(256),
  .DEPTH(4),
  .ADDR_WIDTH(9),
  .GRACE_PERIOD(3)
)
fifo_w_PE_8_9_V_V_U
(
  .clk(ap_clk),
  .reset(ap_rst_n_inv),
  .if_read_ce(1'b1),
  .if_write_ce(1'b1),
  .if_din(PE_wrapper254_U0_fifo_w_out_V_V_din),
  .if_full_n(fifo_w_PE_8_9_V_V_full_n),
  .if_write(PE_wrapper254_U0_fifo_w_out_V_V_write),
  .if_dout(fifo_w_PE_8_9_V_V_dout),
  .if_empty_n(fifo_w_PE_8_9_V_V_empty_n),
  .if_read(PE_wrapper255_U0_fifo_w_in_V_V_read)
);

(* keep_hierarchy = "yes" *)
fifo_almost_full
#(
  .DATA_WIDTH(64),
  .DEPTH(4),
  .ADDR_WIDTH(7),
  .GRACE_PERIOD(3)
)
fifo_cout_drain_cout_drain_IO_L1_out_10_6_V_V_U
(
  .clk(ap_clk),
  .reset(ap_rst_n_inv),
  .if_read_ce(1'b1),
  .if_write_ce(1'b1),
  .if_din(cout_drain_IO_L1_out_wrapper536_U0_fifo_cout_drain_out_V_V_din),
  .if_full_n(fifo_cout_drain_cout_drain_IO_L1_out_10_6_V_V_full_n),
  .if_write(cout_drain_IO_L1_out_wrapper536_U0_fifo_cout_drain_out_V_V_write),
  .if_dout(fifo_cout_drain_cout_drain_IO_L1_out_10_6_V_V_dout),
  .if_empty_n(fifo_cout_drain_cout_drain_IO_L1_out_10_6_V_V_empty_n),
  .if_read(cout_drain_IO_L1_out_wrapper537_U0_fifo_cout_drain_in_V_V_read)
);

(* keep_hierarchy = "yes" *)
fifo_almost_full
#(
  .DATA_WIDTH(256),
  .DEPTH(5),
  .ADDR_WIDTH(9),
  .GRACE_PERIOD(5)
)
fifo_w_PE_2_9_V_V_U
(
  .clk(ap_clk),
  .reset(ap_rst_n_inv),
  .if_read_ce(1'b1),
  .if_write_ce(1'b1),
  .if_din(PE_wrapper182_U0_fifo_w_out_V_V_din),
  .if_full_n(fifo_w_PE_2_9_V_V_full_n),
  .if_write(PE_wrapper182_U0_fifo_w_out_V_V_write),
  .if_dout(fifo_w_PE_2_9_V_V_dout),
  .if_empty_n(fifo_w_PE_2_9_V_V_empty_n),
  .if_read(PE_wrapper183_U0_fifo_w_in_V_V_read)
);

(* keep_hierarchy = "yes" *)
fifo_almost_full
#(
  .DATA_WIDTH(64),
  .DEPTH(5),
  .ADDR_WIDTH(7),
  .GRACE_PERIOD(5)
)
fifo_cout_drain_cout_drain_IO_L1_out_10_8_V_V_U
(
  .clk(ap_clk),
  .reset(ap_rst_n_inv),
  .if_read_ce(1'b1),
  .if_write_ce(1'b1),
  .if_din(cout_drain_IO_L1_out_wrapper534_U0_fifo_cout_drain_out_V_V_din),
  .if_full_n(fifo_cout_drain_cout_drain_IO_L1_out_10_8_V_V_full_n),
  .if_write(cout_drain_IO_L1_out_wrapper534_U0_fifo_cout_drain_out_V_V_write),
  .if_dout(fifo_cout_drain_cout_drain_IO_L1_out_10_8_V_V_dout),
  .if_empty_n(fifo_cout_drain_cout_drain_IO_L1_out_10_8_V_V_empty_n),
  .if_read(cout_drain_IO_L1_out_wrapper535_U0_fifo_cout_drain_in_V_V_read)
);

(* keep_hierarchy = "yes" *)
fifo_almost_full
#(
  .DATA_WIDTH(64),
  .DEPTH(6),
  .ADDR_WIDTH(7),
  .GRACE_PERIOD(7)
)
fifo_cout_drain_cout_drain_IO_L3_out_serialize_V_V_U
(
  .clk(ap_clk),
  .reset(ap_rst_n_inv),
  .if_read_ce(1'b1),
  .if_write_ce(1'b1),
  .if_din(cout_drain_IO_L3_out_U0_fifo_cout_drain_out_V_V_din),
  .if_full_n(fifo_cout_drain_cout_drain_IO_L3_out_serialize_V_V_full_n),
  .if_write(cout_drain_IO_L3_out_U0_fifo_cout_drain_out_V_V_write),
  .if_dout(fifo_cout_drain_cout_drain_IO_L3_out_serialize_V_V_dout),
  .if_empty_n(fifo_cout_drain_cout_drain_IO_L3_out_serialize_V_V_empty_n),
  .if_read(cout_drain_IO_L3_out_serialize_U0_fifo_cout_drain_local_in_V_V_read)
);

(* keep_hierarchy = "yes" *)
fifo_almost_full
#(
  .DATA_WIDTH(256),
  .DEPTH(4),
  .ADDR_WIDTH(9),
  .GRACE_PERIOD(3)
)
fifo_w_PE_5_12_V_V_U
(
  .clk(ap_clk),
  .reset(ap_rst_n_inv),
  .if_read_ce(1'b1),
  .if_write_ce(1'b1),
  .if_din(PE_wrapper221_U0_fifo_w_out_V_V_din),
  .if_full_n(fifo_w_PE_5_12_V_V_full_n),
  .if_write(PE_wrapper221_U0_fifo_w_out_V_V_write),
  .if_dout(fifo_w_PE_5_12_V_V_dout),
  .if_empty_n(fifo_w_PE_5_12_V_V_empty_n),
  .if_read(w_PE_dummy_in357_U0_fifo_w_in_V_V_read)
);

(* keep_hierarchy = "yes" *)
fifo_almost_full
#(
  .DATA_WIDTH(32),
  .DEPTH(53),
  .ADDR_WIDTH(6),
  .GRACE_PERIOD(5)
)
fifo_cout_drain_PE_3_11_V_U
(
  .clk(ap_clk),
  .reset(ap_rst_n_inv),
  .if_read_ce(1'b1),
  .if_write_ce(1'b1),
  .if_din(PE_wrapper197_U0_fifo_cout_drain_out_V_din),
  .if_full_n(fifo_cout_drain_PE_3_11_V_full_n),
  .if_write(PE_wrapper197_U0_fifo_cout_drain_out_V_write),
  .if_dout(fifo_cout_drain_PE_3_11_V_dout),
  .if_empty_n(fifo_cout_drain_PE_3_11_V_empty_n),
  .if_read(cout_drain_IO_L1_out_wrapper554_U0_fifo_cout_drain_local_in_V_read)
);

(* keep_hierarchy = "yes" *)
fifo_almost_full
#(
  .DATA_WIDTH(64),
  .DEPTH(4),
  .ADDR_WIDTH(7),
  .GRACE_PERIOD(3)
)
fifo_cout_drain_cout_drain_IO_L1_out_11_4_V_V_U
(
  .clk(ap_clk),
  .reset(ap_rst_n_inv),
  .if_read_ce(1'b1),
  .if_write_ce(1'b1),
  .if_din(cout_drain_IO_L1_out_wrapper553_U0_fifo_cout_drain_out_V_V_din),
  .if_full_n(fifo_cout_drain_cout_drain_IO_L1_out_11_4_V_V_full_n),
  .if_write(cout_drain_IO_L1_out_wrapper553_U0_fifo_cout_drain_out_V_V_write),
  .if_dout(fifo_cout_drain_cout_drain_IO_L1_out_11_4_V_V_dout),
  .if_empty_n(fifo_cout_drain_cout_drain_IO_L1_out_11_4_V_V_empty_n),
  .if_read(cout_drain_IO_L1_out_wrapper554_U0_fifo_cout_drain_in_V_V_read)
);

// pipeline ap_start
initial begin
  ap_start_p1 = 1'b0;
  ap_start_p2 = 1'b0;
  ap_start_pipe = 1'b0;
end
always @ (posedge ap_clk) begin
  ap_start_p1 <= ap_start;
  ap_start_p2 <= ap_start_p1;
  ap_start_pipe <= ap_start_p2;
end
// pipeline ap_done
always @ (posedge ap_clk) begin
  w_PE_dummy_in357_U0_ap_done_p1 <= w_PE_dummy_in357_U0_ap_done;
  w_PE_dummy_in357_U0_ap_done_p2 <= w_PE_dummy_in357_U0_ap_done_p1;
  w_PE_dummy_in357_U0_ap_done_pipe <= w_PE_dummy_in357_U0_ap_done_p2;
end
always @ (posedge ap_clk) begin
  cout_drain_IO_L3_out_serialize_U0_ap_done_p1 <= cout_drain_IO_L3_out_serialize_U0_ap_done;
  cout_drain_IO_L3_out_serialize_U0_ap_done_p2 <= cout_drain_IO_L3_out_serialize_U0_ap_done_p1;
  cout_drain_IO_L3_out_serialize_U0_ap_done_pipe <= cout_drain_IO_L3_out_serialize_U0_ap_done_p2;
end
(* dont_touch = "yes" *) reg ap_done_reg_;
always @ (posedge ap_clk) begin
  ap_done_reg_ <= w_PE_dummy_in357_U0_ap_done_backup&cout_drain_IO_L3_out_serialize_U0_ap_done_backup;
end
assign ap_done = ap_done_reg_;
// backup ap_done
always @ (posedge ap_clk) begin
  if (ap_done_reg_) begin
    w_PE_dummy_in357_U0_ap_done_backup <= w_PE_dummy_in357_U0_ap_done_pipe;
  end
  else begin
    w_PE_dummy_in357_U0_ap_done_backup <= w_PE_dummy_in357_U0_ap_done_backup | w_PE_dummy_in357_U0_ap_done_pipe;
  end
end
always @ (posedge ap_clk) begin
  if (ap_done_reg_) begin
    cout_drain_IO_L3_out_serialize_U0_ap_done_backup <= cout_drain_IO_L3_out_serialize_U0_ap_done_pipe;
  end
  else begin
    cout_drain_IO_L3_out_serialize_U0_ap_done_backup <= cout_drain_IO_L3_out_serialize_U0_ap_done_backup | cout_drain_IO_L3_out_serialize_U0_ap_done_pipe;
  end
end
assign ap_ready = ap_done;
assign ap_idle = ap_done;
// pipeline ap_start
initial begin
  ap_rst_p1 = 1'b0;
  ap_rst_p2 = 1'b0;
  ap_rst_pipe = 1'b0;
  ap_rst_n_p1 = 1'b0;
  ap_rst_n_p2 = 1'b0;
  ap_rst_n_pipe = 1'b0;
end
always @ (posedge ap_clk) begin
  ap_rst_p1 <= ~ap_rst_n;
  ap_rst_p2 <= ap_rst_p1;
  ap_rst_pipe <= ap_rst_p2;
  ap_rst_n_p1 <= ap_rst_n;
  ap_rst_n_p2 <= ap_rst_n_p1;
  ap_rst_n_pipe <= ap_rst_n_p2;
end
endmodule

// first-word fall-through (FWFT) FIFO
// if its capacity > THRESHOLD bits, it uses block RAM, otherwise it will uses
// shift register LUT
module fifo_almost_full #(
  parameter DATA_WIDTH = 32,
  parameter ADDR_WIDTH = 5,
  parameter DEPTH      = 32,
  parameter THRESHOLD  = 18432,
  parameter GRACE_PERIOD = 2
) (
  input wire clk,
  input wire reset,
  // write
  output wire                  if_full_n,
  input  wire                  if_write_ce,
  input  wire                  if_write,
  input  wire [DATA_WIDTH-1:0] if_din,
  // read
  output wire                  if_empty_n,
  input  wire                  if_read_ce,
  input  wire                  if_read,
  output wire [DATA_WIDTH-1:0] if_dout
);
  parameter REAL_DEPTH = GRACE_PERIOD + DEPTH + 4;
  parameter REAL_ADDR_WIDTH  = $clog2(REAL_DEPTH);
generate
  if (DATA_WIDTH * DEPTH > THRESHOLD) begin : bram
    fifo_bram_almost_full #(
      .DATA_WIDTH(DATA_WIDTH),
      .ADDR_WIDTH(REAL_ADDR_WIDTH),
      .DEPTH     (REAL_DEPTH),
      .GRACE_PERIOD(GRACE_PERIOD) /*********/
    ) unit (
      .clk  (clk),
      .reset(reset),
      .if_full_n  (if_full_n),
      .if_write_ce(if_write_ce),
      .if_write   (if_write),
      .if_din     (if_din),
      .if_empty_n(if_empty_n),
      .if_read_ce(if_read_ce),
      .if_read   (if_read),
      .if_dout   (if_dout)
    );
  end else begin : srl
    fifo_srl_almost_full #(
      .DATA_WIDTH(DATA_WIDTH),
      .ADDR_WIDTH(REAL_ADDR_WIDTH),
      .DEPTH     (REAL_DEPTH),
      .GRACE_PERIOD(GRACE_PERIOD) /*********/
    ) unit (
      .clk  (clk),
      .reset(reset),
      .if_full_n  (if_full_n),
      .if_write_ce(if_write_ce),
      .if_write   (if_write),
      .if_din     (if_din),
      .if_empty_n(if_empty_n),
      .if_read_ce(if_read_ce),
      .if_read   (if_read),
      .if_dout   (if_dout)
    );
  end
endgenerate
endmodule  // fifo
/////////////////////////////////////////////////////////////////
module fifo_srl_almost_full (
    clk,
    reset,
    if_empty_n,
    if_read_ce,
    if_read,
    if_dout,
    if_full_n,
    if_write_ce,
    if_write,
    if_din);
parameter MEM_STYLE   = "shiftreg";
parameter DATA_WIDTH  = 32'd32;
parameter ADDR_WIDTH  = 32'd4;
parameter DEPTH       = 5'd16;
/*******************************************/
parameter GRACE_PERIOD = 2;
/*******************************************/
input clk;
input reset;
output if_empty_n;
input if_read_ce;
input if_read;
output[DATA_WIDTH - 1:0] if_dout;
output if_full_n;
input if_write_ce;
input if_write;
input[DATA_WIDTH - 1:0] if_din;
wire[ADDR_WIDTH - 1:0] shiftReg_addr ;
wire[DATA_WIDTH - 1:0] shiftReg_data, shiftReg_q;
wire                     shiftReg_ce;
reg[ADDR_WIDTH:0] mOutPtr = ~{(ADDR_WIDTH+1){1'b0}};
reg internal_empty_n = 0, internal_full_n = 1;
assign if_empty_n = internal_empty_n;
/*******************************************/
// assign if_full_n = internal_full_n;
wire almost_full = mOutPtr >= DEPTH - 1 - GRACE_PERIOD && mOutPtr != ~{ADDR_WIDTH+1{1'b0}};
assign if_full_n = ~almost_full;
/*******************************************/
assign shiftReg_data = if_din;
assign if_dout = shiftReg_q;
always @ (posedge clk) begin
    if (reset == 1'b1)
    begin
        mOutPtr <= ~{ADDR_WIDTH+1{1'b0}};
        internal_empty_n <= 1'b0;
        internal_full_n <= 1'b1;
    end
    else begin
        if (((if_read & if_read_ce) == 1 & internal_empty_n == 1) && 
            ((if_write & if_write_ce) == 0 | internal_full_n == 0))
        begin
            mOutPtr <= mOutPtr - 5'd1;
            if (mOutPtr == 0)
                internal_empty_n <= 1'b0;
            internal_full_n <= 1'b1;
        end 
        else if (((if_read & if_read_ce) == 0 | internal_empty_n == 0) && 
            ((if_write & if_write_ce) == 1 & internal_full_n == 1))
        begin
            mOutPtr <= mOutPtr + 5'd1;
            internal_empty_n <= 1'b1;
            if (mOutPtr == DEPTH - 5'd2)
                internal_full_n <= 1'b0;
        end 
    end
end
assign shiftReg_addr = mOutPtr[ADDR_WIDTH] == 1'b0 ? mOutPtr[ADDR_WIDTH-1:0]:{ADDR_WIDTH{1'b0}};
assign shiftReg_ce = (if_write & if_write_ce) & internal_full_n;
fifo_srl_almost_full_internal 
#(
    .DATA_WIDTH(DATA_WIDTH),
    .ADDR_WIDTH(ADDR_WIDTH),
    .DEPTH(DEPTH))
U_fifo_w32_d16_A_ram (
    .clk(clk),
    .data(shiftReg_data),
    .ce(shiftReg_ce),
    .a(shiftReg_addr),
    .q(shiftReg_q));
endmodule  
module fifo_srl_almost_full_internal (
    clk,
    data,
    ce,
    a,
    q);
parameter DATA_WIDTH = 32'd32;
parameter ADDR_WIDTH = 32'd4;
parameter DEPTH = 5'd16;
input clk;
input [DATA_WIDTH-1:0] data;
input ce;
input [ADDR_WIDTH-1:0] a;
output [DATA_WIDTH-1:0] q;
reg[DATA_WIDTH-1:0] SRL_SIG [0:DEPTH-1];
integer i;
always @ (posedge clk)
    begin
        if (ce)
        begin
            for (i=0;i<DEPTH-1;i=i+1)
                SRL_SIG[i+1] <= SRL_SIG[i];
            SRL_SIG[0] <= data;
        end
    end
assign q = SRL_SIG[a];
endmodule
///////////////////////////////////////////////////////////
// first-word fall-through (FWFT) FIFO using block RAM or URAM (let Vivado choose)
// based on HLS generated code
module fifo_bram_almost_full #(
  parameter MEM_STYLE  = "auto",
  parameter DATA_WIDTH = 32,
  parameter ADDR_WIDTH = 5,
  parameter DEPTH      = 32,
  parameter GRACE_PERIOD = 2
) (
  input wire clk,
  input wire reset,
  // write
  output wire                  if_full_n,
  input  wire                  if_write_ce,
  input  wire                  if_write,
  input  wire [DATA_WIDTH-1:0] if_din,
  // read
  output wire                  if_empty_n,
  input  wire                  if_read_ce,
  input  wire                  if_read,
  output wire [DATA_WIDTH-1:0] if_dout
);
(* ram_style = MEM_STYLE *)
reg  [DATA_WIDTH-1:0] mem[0:DEPTH-1];
reg  [DATA_WIDTH-1:0] q_buf;
reg  [ADDR_WIDTH-1:0] waddr;
reg  [ADDR_WIDTH-1:0] raddr;
wire [ADDR_WIDTH-1:0] wnext;
wire [ADDR_WIDTH-1:0] rnext;
wire                  push;
wire                  pop;
reg  [ADDR_WIDTH-1:0] used;
reg                   full_n;
reg                   empty_n;
reg  [DATA_WIDTH-1:0] q_tmp;
reg                   show_ahead;
reg  [DATA_WIDTH-1:0] dout_buf;
reg                   dout_valid;
localparam DepthM1 = DEPTH[ADDR_WIDTH-1:0] - 1'd1;
/**************************************/
wire almost_full = (used >= DEPTH - 1 - GRACE_PERIOD);
//assign if_full_n  = full_n;
assign if_full_n  = ~almost_full;
/**************************************/
assign if_empty_n = dout_valid;
assign if_dout    = dout_buf;
assign push       = full_n & if_write_ce & if_write;
assign pop        = empty_n & if_read_ce & (~dout_valid | if_read);
assign wnext      = !push              ? waddr              :
                    (waddr == DepthM1) ? {ADDR_WIDTH{1'b0}} : waddr + 1'd1;
assign rnext      = !pop               ? raddr              :
                    (raddr == DepthM1) ? {ADDR_WIDTH{1'b0}} : raddr + 1'd1;
// waddr
always @(posedge clk) begin
  if (reset)
    waddr <= {ADDR_WIDTH{1'b0}};
  else
    waddr <= wnext;
end
// raddr
always @(posedge clk) begin
  if (reset)
    raddr <= {ADDR_WIDTH{1'b0}};
  else
    raddr <= rnext;
end
// used
always @(posedge clk) begin
  if (reset)
    used <= {ADDR_WIDTH{1'b0}};
  else if (push && !pop)
    used <= used + 1'b1;
  else if (!push && pop)
    used <= used - 1'b1;
end
// full_n
always @(posedge clk) begin
  if (reset)
    full_n <= 1'b1;
  else if (push && !pop)
    full_n <= (used != DepthM1);
  else if (!push && pop)
    full_n <= 1'b1;
end
// empty_n
always @(posedge clk) begin
  if (reset)
    empty_n <= 1'b0;
  else if (push && !pop)
    empty_n <= 1'b1;
  else if (!push && pop)
    empty_n <= (used != {{(ADDR_WIDTH-1){1'b0}},1'b1});
end
// mem
always @(posedge clk) begin
  if (push)
    mem[waddr] <= if_din;
end
// q_buf
always @(posedge clk) begin
  q_buf <= mem[rnext];
end
// q_tmp
always @(posedge clk) begin
  if (reset)
    q_tmp <= {DATA_WIDTH{1'b0}};
  else if (push)
    q_tmp <= if_din;
end
// show_ahead
always @(posedge clk) begin
  if (reset)
    show_ahead <= 1'b0;
  else if (push && used == {{(ADDR_WIDTH-1){1'b0}},pop})
    show_ahead <= 1'b1;
  else
    show_ahead <= 1'b0;
end
// dout_buf
always @(posedge clk) begin
  if (reset)
    dout_buf <= {DATA_WIDTH{1'b0}};
  else if (pop)
    dout_buf <= show_ahead? q_tmp : q_buf;
end
// dout_valid
always @(posedge clk) begin
  if (reset)
    dout_valid <= 1'b0;
  else if (pop)
    dout_valid <= 1'b1;
  else if (if_read_ce & if_read)
    dout_valid <= 1'b0;
end
endmodule  // fifo_bram

