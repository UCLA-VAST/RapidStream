

`timescale 1 ns / 1 ps


module CR_X2Y6_To_CR_X3Y7_ctrl (
  input [31:0] PE_wrapper310_U0_fifo_cout_drain_out_V_din_pass_0,
  output [31:0] PE_wrapper310_U0_fifo_cout_drain_out_V_din_pass_1,
  output fifo_cout_drain_PE_13_4_V_full_n_pass_0,
  input fifo_cout_drain_PE_13_4_V_full_n_pass_1,
  input PE_wrapper310_U0_fifo_cout_drain_out_V_write_pass_0,
  output PE_wrapper310_U0_fifo_cout_drain_out_V_write_pass_1,
  input [31:0] PE_wrapper308_U0_fifo_cout_drain_out_V_din_pass_0,
  output [31:0] PE_wrapper308_U0_fifo_cout_drain_out_V_din_pass_1,
  output fifo_cout_drain_PE_13_2_V_full_n_pass_0,
  input fifo_cout_drain_PE_13_2_V_full_n_pass_1,
  input PE_wrapper308_U0_fifo_cout_drain_out_V_write_pass_0,
  output PE_wrapper308_U0_fifo_cout_drain_out_V_write_pass_1,
  input [255:0] PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0,
  output [255:0] PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_1,
  output fifo_cin_PE_8_4_V_V_full_n_pass_0,
  input fifo_cin_PE_8_4_V_V_full_n_pass_1,
  input PE_wrapper238_U0_fifo_cin_out_V_V_write_pass_0,
  output PE_wrapper238_U0_fifo_cin_out_V_V_write_pass_1,
  input [255:0] PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0,
  output [255:0] PE_wrapper297_U0_fifo_w_out_V_V_din_pass_1,
  output fifo_w_PE_12_4_V_V_full_n_pass_0,
  input fifo_w_PE_12_4_V_V_full_n_pass_1,
  input PE_wrapper297_U0_fifo_w_out_V_V_write_pass_0,
  output PE_wrapper297_U0_fifo_w_out_V_V_write_pass_1,
  input [255:0] PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0,
  output [255:0] PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_1,
  output fifo_cin_PE_14_4_V_V_full_n_pass_0,
  input fifo_cin_PE_14_4_V_V_full_n_pass_1,
  input PE_wrapper310_U0_fifo_cin_out_V_V_write_pass_0,
  output PE_wrapper310_U0_fifo_cin_out_V_V_write_pass_1,
  input [255:0] PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0,
  output [255:0] PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_1,
  output fifo_cin_PE_14_1_V_V_full_n_pass_0,
  input fifo_cin_PE_14_1_V_V_full_n_pass_1,
  input PE_wrapper307_U0_fifo_cin_out_V_V_write_pass_0,
  output PE_wrapper307_U0_fifo_cin_out_V_V_write_pass_1,
  input [255:0] PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0,
  output [255:0] PE_wrapper250_U0_fifo_w_out_V_V_din_pass_1,
  output fifo_w_PE_8_5_V_V_full_n_pass_0,
  input fifo_w_PE_8_5_V_V_full_n_pass_1,
  input PE_wrapper250_U0_fifo_w_out_V_V_write_pass_0,
  output PE_wrapper250_U0_fifo_w_out_V_V_write_pass_1,
  input [255:0] PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0,
  output [255:0] PE_wrapper238_U0_fifo_w_out_V_V_din_pass_1,
  output fifo_w_PE_7_5_V_V_full_n_pass_0,
  input fifo_w_PE_7_5_V_V_full_n_pass_1,
  input PE_wrapper238_U0_fifo_w_out_V_V_write_pass_0,
  output PE_wrapper238_U0_fifo_w_out_V_V_write_pass_1,
  output [31:0] PE_wrapper320_U0_fifo_cout_drain_out_V_din_pass_0,
  input fifo_cout_drain_PE_14_2_V_full_n_pass_0,
  output PE_wrapper320_U0_fifo_cout_drain_out_V_write_pass_0,
  input [63:0] cout_drain_IO_L1_out_wrapper433_U0_fifo_cout_drain_out_V_V_din_pass_0,
  output fifo_cout_drain_cout_drain_IO_L1_out_4_13_V_V_full_n_pass_0,
  input cout_drain_IO_L1_out_wrapper433_U0_fifo_cout_drain_out_V_V_write_pass_0,
  input [255:0] PE_wrapper309_U0_fifo_cin_out_V_V_din_pass_1,
  output fifo_cin_PE_14_3_V_V_full_n_pass_1,
  input PE_wrapper309_U0_fifo_cin_out_V_V_write_pass_1,
  output [63:0] cout_drain_IO_L1_out_wrapper402_U0_fifo_cout_drain_out_V_V_din_pass_0,
  input fifo_cout_drain_cout_drain_IO_L1_out_2_12_V_V_full_n_pass_0,
  output cout_drain_IO_L1_out_wrapper402_U0_fifo_cout_drain_out_V_V_write_pass_0,
  output [255:0] w_IO_L2_in149_U0_fifo_w_out_V_V_din_pass_0,
  input fifo_w_w_IO_L2_in_15_V_V_full_n_pass_0,
  output w_IO_L2_in149_U0_fifo_w_out_V_V_write_pass_0,
  output [31:0] PE_wrapper286_U0_fifo_cout_drain_out_V_din_pass_0,
  input fifo_cout_drain_PE_11_4_V_full_n_pass_0,
  output PE_wrapper286_U0_fifo_cout_drain_out_V_write_pass_0,
  input [255:0] PE_wrapper214_U0_fifo_cin_out_V_V_din_pass_1,
  output fifo_cin_PE_6_4_V_V_full_n_pass_1,
  input PE_wrapper214_U0_fifo_cin_out_V_V_write_pass_1,
  output [63:0] cout_drain_IO_L1_out_wrapper432_U0_fifo_cout_drain_out_V_V_din_pass_0,
  input fifo_cout_drain_cout_drain_IO_L1_out_4_14_V_V_full_n_pass_0,
  output cout_drain_IO_L1_out_wrapper432_U0_fifo_cout_drain_out_V_V_write_pass_0,
  output [255:0] PE_wrapper318_U0_fifo_w_out_V_V_din_pass_0,
  input fifo_w_PE_14_1_V_V_full_n_pass_0,
  output PE_wrapper318_U0_fifo_w_out_V_V_write_pass_0,
  output [31:0] PE_wrapper226_U0_fifo_cout_drain_out_V_din_pass_0,
  input fifo_cout_drain_PE_6_4_V_full_n_pass_0,
  output PE_wrapper226_U0_fifo_cout_drain_out_V_write_pass_0,
  output [255:0] PE_wrapper286_U0_fifo_cin_out_V_V_din_pass_0,
  input fifo_cin_PE_12_4_V_V_full_n_pass_0,
  output PE_wrapper286_U0_fifo_cin_out_V_V_write_pass_0,
  input [255:0] w_IO_L2_in148_U0_fifo_w_out_V_V_din_pass_0,
  output fifo_w_w_IO_L2_in_14_V_V_full_n_pass_0,
  input w_IO_L2_in148_U0_fifo_w_out_V_V_write_pass_0,
  output [255:0] PE_wrapper320_U0_fifo_cin_out_V_V_din_pass_0,
  input fifo_cin_PE_15_2_V_V_full_n_pass_0,
  output PE_wrapper320_U0_fifo_cin_out_V_V_write_pass_0,
  input [63:0] cout_drain_IO_L1_out_wrapper418_U0_fifo_cout_drain_out_V_V_din_pass_1,
  output fifo_cout_drain_cout_drain_IO_L1_out_3_12_V_V_full_n_pass_1,
  input cout_drain_IO_L1_out_wrapper418_U0_fifo_cout_drain_out_V_V_write_pass_1,
  input [255:0] PE_wrapper225_U0_fifo_w_out_V_V_din_pass_1,
  output fifo_w_PE_6_4_V_V_full_n_pass_1,
  input PE_wrapper225_U0_fifo_w_out_V_V_write_pass_1,
  output [63:0] cout_drain_IO_L1_out_wrapper416_U0_fifo_cout_drain_out_V_V_din_pass_0,
  input fifo_cout_drain_cout_drain_IO_L1_out_3_14_V_V_full_n_pass_0,
  output cout_drain_IO_L1_out_wrapper416_U0_fifo_cout_drain_out_V_V_write_pass_0,
  output [255:0] PE_wrapper330_U0_fifo_cin_out_V_V_din_pass_0,
  input fifo_cin_PE_16_0_V_V_full_n_pass_0,
  output PE_wrapper330_U0_fifo_cin_out_V_V_write_pass_0,
  output [255:0] PE_wrapper330_U0_fifo_w_out_V_V_din_pass_0,
  input fifo_w_PE_15_1_V_V_full_n_pass_0,
  output PE_wrapper330_U0_fifo_w_out_V_V_write_pass_0,
  input [255:0] PE_wrapper285_U0_fifo_w_out_V_V_din_pass_1,
  output fifo_w_PE_11_4_V_V_full_n_pass_1,
  input PE_wrapper285_U0_fifo_w_out_V_V_write_pass_1,
  output [63:0] cout_drain_IO_L1_out_wrapper419_U0_fifo_cout_drain_out_V_V_din_pass_0,
  input fifo_cout_drain_cout_drain_IO_L1_out_3_11_V_V_full_n_pass_0,
  output cout_drain_IO_L1_out_wrapper419_U0_fifo_cout_drain_out_V_V_write_pass_0,
  input [255:0] w_IO_L2_in_boundary_U0_fifo_w_local_out_V_V_din_pass_0,
  output fifo_w_PE_15_0_V_V_full_n_pass_0,
  input w_IO_L2_in_boundary_U0_fifo_w_local_out_V_V_write_pass_0,
  input [255:0] PE_wrapper273_U0_fifo_w_out_V_V_din_pass_0,
  output fifo_w_PE_10_4_V_V_full_n_pass_0,
  input PE_wrapper273_U0_fifo_w_out_V_V_write_pass_0,
  output [255:0] PE_wrapper286_U0_fifo_w_out_V_V_din_pass_0,
  input fifo_w_PE_11_5_V_V_full_n_pass_0,
  output PE_wrapper286_U0_fifo_w_out_V_V_write_pass_0,
  input [63:0] cout_drain_IO_L1_out_boundary_wrapper383_U0_fifo_cout_drain_out_V_V_din_pass_0,
  output fifo_cout_drain_cout_drain_IO_L1_out_1_15_V_V_full_n_pass_0,
  input cout_drain_IO_L1_out_boundary_wrapper383_U0_fifo_cout_drain_out_V_V_write_pass_0,
  output [31:0] PE_wrapper330_U0_fifo_cout_drain_out_V_din_pass_0,
  input fifo_cout_drain_PE_15_0_V_full_n_pass_0,
  output PE_wrapper330_U0_fifo_cout_drain_out_V_write_pass_0,
  input [255:0] PE_wrapper306_U0_fifo_cin_out_V_V_din_pass_1,
  output fifo_cin_PE_14_0_V_V_full_n_pass_1,
  input PE_wrapper306_U0_fifo_cin_out_V_V_write_pass_1,
  output [255:0] PE_wrapper321_U0_fifo_cin_out_V_V_din_pass_0,
  input fifo_cin_PE_15_3_V_V_full_n_pass_0,
  output PE_wrapper321_U0_fifo_cin_out_V_V_write_pass_0,
  input [31:0] PE_wrapper285_U0_fifo_cout_drain_out_V_din_pass_1,
  output fifo_cout_drain_PE_11_3_V_full_n_pass_1,
  input PE_wrapper285_U0_fifo_cout_drain_out_V_write_pass_1,
  input [255:0] PE_wrapper319_U0_fifo_w_out_V_V_din_pass_0,
  output fifo_w_PE_14_2_V_V_full_n_pass_0,
  input PE_wrapper319_U0_fifo_w_out_V_V_write_pass_0,
  output [255:0] PE_wrapper226_U0_fifo_w_out_V_V_din_pass_0,
  input fifo_w_PE_6_5_V_V_full_n_pass_0,
  output PE_wrapper226_U0_fifo_w_out_V_V_write_pass_0,
  input [255:0] PE_wrapper308_U0_fifo_cin_out_V_V_din_pass_0,
  output fifo_cin_PE_14_2_V_V_full_n_pass_0,
  input PE_wrapper308_U0_fifo_cin_out_V_V_write_pass_0,
  output [63:0] cout_drain_IO_L1_out_wrapper384_U0_fifo_cout_drain_out_V_V_din_pass_0,
  input fifo_cout_drain_cout_drain_IO_L1_out_1_14_V_V_full_n_pass_0,
  output cout_drain_IO_L1_out_wrapper384_U0_fifo_cout_drain_out_V_V_write_pass_0,
  input [31:0] PE_wrapper319_U0_fifo_cout_drain_out_V_din_pass_0,
  output fifo_cout_drain_PE_14_1_V_full_n_pass_0,
  input PE_wrapper319_U0_fifo_cout_drain_out_V_write_pass_0,
  input [31:0] PE_wrapper334_U0_fifo_cout_drain_out_V_din_pass_0,
  output fifo_cout_drain_PE_15_4_V_full_n_pass_0,
  input PE_wrapper334_U0_fifo_cout_drain_out_V_write_pass_0,
  input [63:0] cout_drain_IO_L1_out_boundary_wrapper415_U0_fifo_cout_drain_out_V_V_din_pass_0,
  output fifo_cout_drain_cout_drain_IO_L1_out_3_15_V_V_full_n_pass_0,
  input cout_drain_IO_L1_out_boundary_wrapper415_U0_fifo_cout_drain_out_V_V_write_pass_0,
  output [255:0] PE_wrapper274_U0_fifo_w_out_V_V_din_pass_0,
  input fifo_w_PE_10_5_V_V_full_n_pass_0,
  output PE_wrapper274_U0_fifo_w_out_V_V_write_pass_0,
  input [255:0] PE_wrapper262_U0_fifo_cin_out_V_V_din_pass_1,
  output fifo_cin_PE_10_4_V_V_full_n_pass_1,
  input PE_wrapper262_U0_fifo_cin_out_V_V_write_pass_1,
  output [255:0] PE_wrapper226_U0_fifo_cin_out_V_V_din_pass_0,
  input fifo_cin_PE_7_4_V_V_full_n_pass_0,
  output PE_wrapper226_U0_fifo_cin_out_V_V_write_pass_0,
  output [31:0] PE_wrapper318_U0_fifo_cout_drain_out_V_din_pass_0,
  input fifo_cout_drain_PE_14_0_V_full_n_pass_0,
  output PE_wrapper318_U0_fifo_cout_drain_out_V_write_pass_0,
  output [31:0] PE_wrapper274_U0_fifo_cout_drain_out_V_din_pass_0,
  input fifo_cout_drain_PE_10_4_V_full_n_pass_0,
  output PE_wrapper274_U0_fifo_cout_drain_out_V_write_pass_0,
  input [31:0] PE_wrapper296_U0_fifo_cout_drain_out_V_din_pass_1,
  output fifo_cout_drain_PE_12_2_V_full_n_pass_1,
  input PE_wrapper296_U0_fifo_cout_drain_out_V_write_pass_1,
  output [255:0] PE_wrapper321_U0_fifo_w_out_V_V_din_pass_0,
  input fifo_w_PE_14_4_V_V_full_n_pass_0,
  output PE_wrapper321_U0_fifo_w_out_V_V_write_pass_0,
  input [31:0] PE_wrapper322_U0_fifo_cout_drain_out_V_din_pass_0,
  output fifo_cout_drain_PE_14_4_V_full_n_pass_0,
  input PE_wrapper322_U0_fifo_cout_drain_out_V_write_pass_0,
  input [63:0] cout_drain_IO_L1_out_wrapper401_U0_fifo_cout_drain_out_V_V_din_pass_0,
  output fifo_cout_drain_cout_drain_IO_L1_out_2_13_V_V_full_n_pass_0,
  input cout_drain_IO_L1_out_wrapper401_U0_fifo_cout_drain_out_V_V_write_pass_0,
  output [63:0] cout_drain_IO_L1_out_wrapper434_U0_fifo_cout_drain_out_V_V_din_pass_0,
  input fifo_cout_drain_cout_drain_IO_L1_out_4_12_V_V_full_n_pass_0,
  output cout_drain_IO_L1_out_wrapper434_U0_fifo_cout_drain_out_V_V_write_pass_0,
  input [31:0] PE_wrapper298_U0_fifo_cout_drain_out_V_din_pass_0,
  output fifo_cout_drain_PE_12_4_V_full_n_pass_0,
  input PE_wrapper298_U0_fifo_cout_drain_out_V_write_pass_0,
  input ap_clk,
  input ap_start_Boundary_X2Y6_To_X4Y6,
  input ap_rst_n_Boundary_X2Y6_To_X4Y6,
  output ap_done_Boundary_X2Y6_To_X4Y6,
  output ap_start_Boundary_X2Y8_To_X4Y8,
  output ap_rst_n_Boundary_X2Y8_To_X4Y8,
  input ap_done_Boundary_X2Y8_To_X4Y8
);
wire ap_start;
wire ap_rst_n;
wire ap_done;
wire ap_idle;
wire ap_ready;
wire ap_continue = 1;
(* keep = "true" *) reg ap_start_Boundary_X2Y6_To_X4Y6_q;
always @ (posedge ap_clk) ap_start_Boundary_X2Y6_To_X4Y6_q <= ap_start_Boundary_X2Y6_To_X4Y6;
assign ap_start_Boundary_X2Y8_To_X4Y8 = ap_start_Boundary_X2Y6_To_X4Y6_q;
assign ap_start = ap_start_Boundary_X2Y6_To_X4Y6_q;
(* keep = "true" *) reg ap_rst_n_Boundary_X2Y6_To_X4Y6_q;
always @ (posedge ap_clk) ap_rst_n_Boundary_X2Y6_To_X4Y6_q <= ap_rst_n_Boundary_X2Y6_To_X4Y6;
assign ap_rst_n_Boundary_X2Y8_To_X4Y8 = ap_rst_n_Boundary_X2Y6_To_X4Y6_q;
assign ap_rst_n = ap_rst_n_Boundary_X2Y6_To_X4Y6_q;
(* keep = "true" *) reg ap_done_Boundary_X2Y8_To_X4Y8_q;
always @ (posedge ap_clk) begin
  if (!ap_rst_n) ap_done_Boundary_X2Y8_To_X4Y8_q <= 0;
  else ap_done_Boundary_X2Y8_To_X4Y8_q <= ap_done_Boundary_X2Y8_To_X4Y8_q | ap_done_Boundary_X2Y8_To_X4Y8;
end
assign ap_done_Boundary_X2Y6_To_X4Y6 = ap_done_Boundary_X2Y8_To_X4Y8_q & ap_done;


  (* dont_touch = "yes" *) CR_X2Y6_To_CR_X3Y7_routing CR_X2Y6_To_CR_X3Y7_routing_U0 (
    .PE_wrapper310_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper310_U0_fifo_cout_drain_out_V_din_pass_0),
    .PE_wrapper310_U0_fifo_cout_drain_out_V_din_pass_1(PE_wrapper310_U0_fifo_cout_drain_out_V_din_pass_1),
    .fifo_cout_drain_PE_13_4_V_full_n_pass_0(fifo_cout_drain_PE_13_4_V_full_n_pass_0),
    .fifo_cout_drain_PE_13_4_V_full_n_pass_1(fifo_cout_drain_PE_13_4_V_full_n_pass_1),
    .PE_wrapper310_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper310_U0_fifo_cout_drain_out_V_write_pass_0),
    .PE_wrapper310_U0_fifo_cout_drain_out_V_write_pass_1(PE_wrapper310_U0_fifo_cout_drain_out_V_write_pass_1),
    .PE_wrapper308_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper308_U0_fifo_cout_drain_out_V_din_pass_0),
    .PE_wrapper308_U0_fifo_cout_drain_out_V_din_pass_1(PE_wrapper308_U0_fifo_cout_drain_out_V_din_pass_1),
    .fifo_cout_drain_PE_13_2_V_full_n_pass_0(fifo_cout_drain_PE_13_2_V_full_n_pass_0),
    .fifo_cout_drain_PE_13_2_V_full_n_pass_1(fifo_cout_drain_PE_13_2_V_full_n_pass_1),
    .PE_wrapper308_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper308_U0_fifo_cout_drain_out_V_write_pass_0),
    .PE_wrapper308_U0_fifo_cout_drain_out_V_write_pass_1(PE_wrapper308_U0_fifo_cout_drain_out_V_write_pass_1),
    .PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0),
    .PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_1(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_1),
    .fifo_cin_PE_8_4_V_V_full_n_pass_0(fifo_cin_PE_8_4_V_V_full_n_pass_0),
    .fifo_cin_PE_8_4_V_V_full_n_pass_1(fifo_cin_PE_8_4_V_V_full_n_pass_1),
    .PE_wrapper238_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper238_U0_fifo_cin_out_V_V_write_pass_0),
    .PE_wrapper238_U0_fifo_cin_out_V_V_write_pass_1(PE_wrapper238_U0_fifo_cin_out_V_V_write_pass_1),
    .PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0),
    .PE_wrapper297_U0_fifo_w_out_V_V_din_pass_1(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_1),
    .fifo_w_PE_12_4_V_V_full_n_pass_0(fifo_w_PE_12_4_V_V_full_n_pass_0),
    .fifo_w_PE_12_4_V_V_full_n_pass_1(fifo_w_PE_12_4_V_V_full_n_pass_1),
    .PE_wrapper297_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper297_U0_fifo_w_out_V_V_write_pass_0),
    .PE_wrapper297_U0_fifo_w_out_V_V_write_pass_1(PE_wrapper297_U0_fifo_w_out_V_V_write_pass_1),
    .PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0),
    .PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_1(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_1),
    .fifo_cin_PE_14_4_V_V_full_n_pass_0(fifo_cin_PE_14_4_V_V_full_n_pass_0),
    .fifo_cin_PE_14_4_V_V_full_n_pass_1(fifo_cin_PE_14_4_V_V_full_n_pass_1),
    .PE_wrapper310_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper310_U0_fifo_cin_out_V_V_write_pass_0),
    .PE_wrapper310_U0_fifo_cin_out_V_V_write_pass_1(PE_wrapper310_U0_fifo_cin_out_V_V_write_pass_1),
    .PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0),
    .PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_1(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_1),
    .fifo_cin_PE_14_1_V_V_full_n_pass_0(fifo_cin_PE_14_1_V_V_full_n_pass_0),
    .fifo_cin_PE_14_1_V_V_full_n_pass_1(fifo_cin_PE_14_1_V_V_full_n_pass_1),
    .PE_wrapper307_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper307_U0_fifo_cin_out_V_V_write_pass_0),
    .PE_wrapper307_U0_fifo_cin_out_V_V_write_pass_1(PE_wrapper307_U0_fifo_cin_out_V_V_write_pass_1),
    .PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0),
    .PE_wrapper250_U0_fifo_w_out_V_V_din_pass_1(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_1),
    .fifo_w_PE_8_5_V_V_full_n_pass_0(fifo_w_PE_8_5_V_V_full_n_pass_0),
    .fifo_w_PE_8_5_V_V_full_n_pass_1(fifo_w_PE_8_5_V_V_full_n_pass_1),
    .PE_wrapper250_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper250_U0_fifo_w_out_V_V_write_pass_0),
    .PE_wrapper250_U0_fifo_w_out_V_V_write_pass_1(PE_wrapper250_U0_fifo_w_out_V_V_write_pass_1),
    .PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0),
    .PE_wrapper238_U0_fifo_w_out_V_V_din_pass_1(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_1),
    .fifo_w_PE_7_5_V_V_full_n_pass_0(fifo_w_PE_7_5_V_V_full_n_pass_0),
    .fifo_w_PE_7_5_V_V_full_n_pass_1(fifo_w_PE_7_5_V_V_full_n_pass_1),
    .PE_wrapper238_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper238_U0_fifo_w_out_V_V_write_pass_0),
    .PE_wrapper238_U0_fifo_w_out_V_V_write_pass_1(PE_wrapper238_U0_fifo_w_out_V_V_write_pass_1),
    .PE_wrapper320_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper320_U0_fifo_cout_drain_out_V_din_pass_0),
    .fifo_cout_drain_PE_14_2_V_full_n_pass_0(fifo_cout_drain_PE_14_2_V_full_n_pass_0),
    .PE_wrapper320_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper320_U0_fifo_cout_drain_out_V_write_pass_0),
    .cout_drain_IO_L1_out_wrapper433_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper433_U0_fifo_cout_drain_out_V_V_din_pass_0),
    .fifo_cout_drain_cout_drain_IO_L1_out_4_13_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_4_13_V_V_full_n_pass_0),
    .cout_drain_IO_L1_out_wrapper433_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper433_U0_fifo_cout_drain_out_V_V_write_pass_0),
    .PE_wrapper309_U0_fifo_cin_out_V_V_din_pass_1(PE_wrapper309_U0_fifo_cin_out_V_V_din_pass_1),
    .fifo_cin_PE_14_3_V_V_full_n_pass_1(fifo_cin_PE_14_3_V_V_full_n_pass_1),
    .PE_wrapper309_U0_fifo_cin_out_V_V_write_pass_1(PE_wrapper309_U0_fifo_cin_out_V_V_write_pass_1),
    .cout_drain_IO_L1_out_wrapper402_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper402_U0_fifo_cout_drain_out_V_V_din_pass_0),
    .fifo_cout_drain_cout_drain_IO_L1_out_2_12_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_2_12_V_V_full_n_pass_0),
    .cout_drain_IO_L1_out_wrapper402_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper402_U0_fifo_cout_drain_out_V_V_write_pass_0),
    .w_IO_L2_in149_U0_fifo_w_out_V_V_din_pass_0(w_IO_L2_in149_U0_fifo_w_out_V_V_din_pass_0),
    .fifo_w_w_IO_L2_in_15_V_V_full_n_pass_0(fifo_w_w_IO_L2_in_15_V_V_full_n_pass_0),
    .w_IO_L2_in149_U0_fifo_w_out_V_V_write_pass_0(w_IO_L2_in149_U0_fifo_w_out_V_V_write_pass_0),
    .PE_wrapper286_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper286_U0_fifo_cout_drain_out_V_din_pass_0),
    .fifo_cout_drain_PE_11_4_V_full_n_pass_0(fifo_cout_drain_PE_11_4_V_full_n_pass_0),
    .PE_wrapper286_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper286_U0_fifo_cout_drain_out_V_write_pass_0),
    .PE_wrapper214_U0_fifo_cin_out_V_V_din_pass_1(PE_wrapper214_U0_fifo_cin_out_V_V_din_pass_1),
    .fifo_cin_PE_6_4_V_V_full_n_pass_1(fifo_cin_PE_6_4_V_V_full_n_pass_1),
    .PE_wrapper214_U0_fifo_cin_out_V_V_write_pass_1(PE_wrapper214_U0_fifo_cin_out_V_V_write_pass_1),
    .cout_drain_IO_L1_out_wrapper432_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper432_U0_fifo_cout_drain_out_V_V_din_pass_0),
    .fifo_cout_drain_cout_drain_IO_L1_out_4_14_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_4_14_V_V_full_n_pass_0),
    .cout_drain_IO_L1_out_wrapper432_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper432_U0_fifo_cout_drain_out_V_V_write_pass_0),
    .PE_wrapper318_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper318_U0_fifo_w_out_V_V_din_pass_0),
    .fifo_w_PE_14_1_V_V_full_n_pass_0(fifo_w_PE_14_1_V_V_full_n_pass_0),
    .PE_wrapper318_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper318_U0_fifo_w_out_V_V_write_pass_0),
    .PE_wrapper226_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper226_U0_fifo_cout_drain_out_V_din_pass_0),
    .fifo_cout_drain_PE_6_4_V_full_n_pass_0(fifo_cout_drain_PE_6_4_V_full_n_pass_0),
    .PE_wrapper226_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper226_U0_fifo_cout_drain_out_V_write_pass_0),
    .PE_wrapper286_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper286_U0_fifo_cin_out_V_V_din_pass_0),
    .fifo_cin_PE_12_4_V_V_full_n_pass_0(fifo_cin_PE_12_4_V_V_full_n_pass_0),
    .PE_wrapper286_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper286_U0_fifo_cin_out_V_V_write_pass_0),
    .w_IO_L2_in148_U0_fifo_w_out_V_V_din_pass_0(w_IO_L2_in148_U0_fifo_w_out_V_V_din_pass_0),
    .fifo_w_w_IO_L2_in_14_V_V_full_n_pass_0(fifo_w_w_IO_L2_in_14_V_V_full_n_pass_0),
    .w_IO_L2_in148_U0_fifo_w_out_V_V_write_pass_0(w_IO_L2_in148_U0_fifo_w_out_V_V_write_pass_0),
    .PE_wrapper320_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper320_U0_fifo_cin_out_V_V_din_pass_0),
    .fifo_cin_PE_15_2_V_V_full_n_pass_0(fifo_cin_PE_15_2_V_V_full_n_pass_0),
    .PE_wrapper320_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper320_U0_fifo_cin_out_V_V_write_pass_0),
    .cout_drain_IO_L1_out_wrapper418_U0_fifo_cout_drain_out_V_V_din_pass_1(cout_drain_IO_L1_out_wrapper418_U0_fifo_cout_drain_out_V_V_din_pass_1),
    .fifo_cout_drain_cout_drain_IO_L1_out_3_12_V_V_full_n_pass_1(fifo_cout_drain_cout_drain_IO_L1_out_3_12_V_V_full_n_pass_1),
    .cout_drain_IO_L1_out_wrapper418_U0_fifo_cout_drain_out_V_V_write_pass_1(cout_drain_IO_L1_out_wrapper418_U0_fifo_cout_drain_out_V_V_write_pass_1),
    .PE_wrapper225_U0_fifo_w_out_V_V_din_pass_1(PE_wrapper225_U0_fifo_w_out_V_V_din_pass_1),
    .fifo_w_PE_6_4_V_V_full_n_pass_1(fifo_w_PE_6_4_V_V_full_n_pass_1),
    .PE_wrapper225_U0_fifo_w_out_V_V_write_pass_1(PE_wrapper225_U0_fifo_w_out_V_V_write_pass_1),
    .cout_drain_IO_L1_out_wrapper416_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper416_U0_fifo_cout_drain_out_V_V_din_pass_0),
    .fifo_cout_drain_cout_drain_IO_L1_out_3_14_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_3_14_V_V_full_n_pass_0),
    .cout_drain_IO_L1_out_wrapper416_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper416_U0_fifo_cout_drain_out_V_V_write_pass_0),
    .PE_wrapper330_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper330_U0_fifo_cin_out_V_V_din_pass_0),
    .fifo_cin_PE_16_0_V_V_full_n_pass_0(fifo_cin_PE_16_0_V_V_full_n_pass_0),
    .PE_wrapper330_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper330_U0_fifo_cin_out_V_V_write_pass_0),
    .PE_wrapper330_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper330_U0_fifo_w_out_V_V_din_pass_0),
    .fifo_w_PE_15_1_V_V_full_n_pass_0(fifo_w_PE_15_1_V_V_full_n_pass_0),
    .PE_wrapper330_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper330_U0_fifo_w_out_V_V_write_pass_0),
    .PE_wrapper285_U0_fifo_w_out_V_V_din_pass_1(PE_wrapper285_U0_fifo_w_out_V_V_din_pass_1),
    .fifo_w_PE_11_4_V_V_full_n_pass_1(fifo_w_PE_11_4_V_V_full_n_pass_1),
    .PE_wrapper285_U0_fifo_w_out_V_V_write_pass_1(PE_wrapper285_U0_fifo_w_out_V_V_write_pass_1),
    .cout_drain_IO_L1_out_wrapper419_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper419_U0_fifo_cout_drain_out_V_V_din_pass_0),
    .fifo_cout_drain_cout_drain_IO_L1_out_3_11_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_3_11_V_V_full_n_pass_0),
    .cout_drain_IO_L1_out_wrapper419_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper419_U0_fifo_cout_drain_out_V_V_write_pass_0),
    .w_IO_L2_in_boundary_U0_fifo_w_local_out_V_V_din_pass_0(w_IO_L2_in_boundary_U0_fifo_w_local_out_V_V_din_pass_0),
    .fifo_w_PE_15_0_V_V_full_n_pass_0(fifo_w_PE_15_0_V_V_full_n_pass_0),
    .w_IO_L2_in_boundary_U0_fifo_w_local_out_V_V_write_pass_0(w_IO_L2_in_boundary_U0_fifo_w_local_out_V_V_write_pass_0),
    .PE_wrapper273_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper273_U0_fifo_w_out_V_V_din_pass_0),
    .fifo_w_PE_10_4_V_V_full_n_pass_0(fifo_w_PE_10_4_V_V_full_n_pass_0),
    .PE_wrapper273_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper273_U0_fifo_w_out_V_V_write_pass_0),
    .PE_wrapper286_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper286_U0_fifo_w_out_V_V_din_pass_0),
    .fifo_w_PE_11_5_V_V_full_n_pass_0(fifo_w_PE_11_5_V_V_full_n_pass_0),
    .PE_wrapper286_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper286_U0_fifo_w_out_V_V_write_pass_0),
    .cout_drain_IO_L1_out_boundary_wrapper383_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_boundary_wrapper383_U0_fifo_cout_drain_out_V_V_din_pass_0),
    .fifo_cout_drain_cout_drain_IO_L1_out_1_15_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_1_15_V_V_full_n_pass_0),
    .cout_drain_IO_L1_out_boundary_wrapper383_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_boundary_wrapper383_U0_fifo_cout_drain_out_V_V_write_pass_0),
    .PE_wrapper330_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper330_U0_fifo_cout_drain_out_V_din_pass_0),
    .fifo_cout_drain_PE_15_0_V_full_n_pass_0(fifo_cout_drain_PE_15_0_V_full_n_pass_0),
    .PE_wrapper330_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper330_U0_fifo_cout_drain_out_V_write_pass_0),
    .PE_wrapper306_U0_fifo_cin_out_V_V_din_pass_1(PE_wrapper306_U0_fifo_cin_out_V_V_din_pass_1),
    .fifo_cin_PE_14_0_V_V_full_n_pass_1(fifo_cin_PE_14_0_V_V_full_n_pass_1),
    .PE_wrapper306_U0_fifo_cin_out_V_V_write_pass_1(PE_wrapper306_U0_fifo_cin_out_V_V_write_pass_1),
    .PE_wrapper321_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper321_U0_fifo_cin_out_V_V_din_pass_0),
    .fifo_cin_PE_15_3_V_V_full_n_pass_0(fifo_cin_PE_15_3_V_V_full_n_pass_0),
    .PE_wrapper321_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper321_U0_fifo_cin_out_V_V_write_pass_0),
    .PE_wrapper285_U0_fifo_cout_drain_out_V_din_pass_1(PE_wrapper285_U0_fifo_cout_drain_out_V_din_pass_1),
    .fifo_cout_drain_PE_11_3_V_full_n_pass_1(fifo_cout_drain_PE_11_3_V_full_n_pass_1),
    .PE_wrapper285_U0_fifo_cout_drain_out_V_write_pass_1(PE_wrapper285_U0_fifo_cout_drain_out_V_write_pass_1),
    .PE_wrapper319_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper319_U0_fifo_w_out_V_V_din_pass_0),
    .fifo_w_PE_14_2_V_V_full_n_pass_0(fifo_w_PE_14_2_V_V_full_n_pass_0),
    .PE_wrapper319_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper319_U0_fifo_w_out_V_V_write_pass_0),
    .PE_wrapper226_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper226_U0_fifo_w_out_V_V_din_pass_0),
    .fifo_w_PE_6_5_V_V_full_n_pass_0(fifo_w_PE_6_5_V_V_full_n_pass_0),
    .PE_wrapper226_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper226_U0_fifo_w_out_V_V_write_pass_0),
    .PE_wrapper308_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper308_U0_fifo_cin_out_V_V_din_pass_0),
    .fifo_cin_PE_14_2_V_V_full_n_pass_0(fifo_cin_PE_14_2_V_V_full_n_pass_0),
    .PE_wrapper308_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper308_U0_fifo_cin_out_V_V_write_pass_0),
    .cout_drain_IO_L1_out_wrapper384_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper384_U0_fifo_cout_drain_out_V_V_din_pass_0),
    .fifo_cout_drain_cout_drain_IO_L1_out_1_14_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_1_14_V_V_full_n_pass_0),
    .cout_drain_IO_L1_out_wrapper384_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper384_U0_fifo_cout_drain_out_V_V_write_pass_0),
    .PE_wrapper319_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper319_U0_fifo_cout_drain_out_V_din_pass_0),
    .fifo_cout_drain_PE_14_1_V_full_n_pass_0(fifo_cout_drain_PE_14_1_V_full_n_pass_0),
    .PE_wrapper319_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper319_U0_fifo_cout_drain_out_V_write_pass_0),
    .PE_wrapper334_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper334_U0_fifo_cout_drain_out_V_din_pass_0),
    .fifo_cout_drain_PE_15_4_V_full_n_pass_0(fifo_cout_drain_PE_15_4_V_full_n_pass_0),
    .PE_wrapper334_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper334_U0_fifo_cout_drain_out_V_write_pass_0),
    .cout_drain_IO_L1_out_boundary_wrapper415_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_boundary_wrapper415_U0_fifo_cout_drain_out_V_V_din_pass_0),
    .fifo_cout_drain_cout_drain_IO_L1_out_3_15_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_3_15_V_V_full_n_pass_0),
    .cout_drain_IO_L1_out_boundary_wrapper415_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_boundary_wrapper415_U0_fifo_cout_drain_out_V_V_write_pass_0),
    .PE_wrapper274_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper274_U0_fifo_w_out_V_V_din_pass_0),
    .fifo_w_PE_10_5_V_V_full_n_pass_0(fifo_w_PE_10_5_V_V_full_n_pass_0),
    .PE_wrapper274_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper274_U0_fifo_w_out_V_V_write_pass_0),
    .PE_wrapper262_U0_fifo_cin_out_V_V_din_pass_1(PE_wrapper262_U0_fifo_cin_out_V_V_din_pass_1),
    .fifo_cin_PE_10_4_V_V_full_n_pass_1(fifo_cin_PE_10_4_V_V_full_n_pass_1),
    .PE_wrapper262_U0_fifo_cin_out_V_V_write_pass_1(PE_wrapper262_U0_fifo_cin_out_V_V_write_pass_1),
    .PE_wrapper226_U0_fifo_cin_out_V_V_din_pass_0(PE_wrapper226_U0_fifo_cin_out_V_V_din_pass_0),
    .fifo_cin_PE_7_4_V_V_full_n_pass_0(fifo_cin_PE_7_4_V_V_full_n_pass_0),
    .PE_wrapper226_U0_fifo_cin_out_V_V_write_pass_0(PE_wrapper226_U0_fifo_cin_out_V_V_write_pass_0),
    .PE_wrapper318_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper318_U0_fifo_cout_drain_out_V_din_pass_0),
    .fifo_cout_drain_PE_14_0_V_full_n_pass_0(fifo_cout_drain_PE_14_0_V_full_n_pass_0),
    .PE_wrapper318_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper318_U0_fifo_cout_drain_out_V_write_pass_0),
    .PE_wrapper274_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper274_U0_fifo_cout_drain_out_V_din_pass_0),
    .fifo_cout_drain_PE_10_4_V_full_n_pass_0(fifo_cout_drain_PE_10_4_V_full_n_pass_0),
    .PE_wrapper274_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper274_U0_fifo_cout_drain_out_V_write_pass_0),
    .PE_wrapper296_U0_fifo_cout_drain_out_V_din_pass_1(PE_wrapper296_U0_fifo_cout_drain_out_V_din_pass_1),
    .fifo_cout_drain_PE_12_2_V_full_n_pass_1(fifo_cout_drain_PE_12_2_V_full_n_pass_1),
    .PE_wrapper296_U0_fifo_cout_drain_out_V_write_pass_1(PE_wrapper296_U0_fifo_cout_drain_out_V_write_pass_1),
    .PE_wrapper321_U0_fifo_w_out_V_V_din_pass_0(PE_wrapper321_U0_fifo_w_out_V_V_din_pass_0),
    .fifo_w_PE_14_4_V_V_full_n_pass_0(fifo_w_PE_14_4_V_V_full_n_pass_0),
    .PE_wrapper321_U0_fifo_w_out_V_V_write_pass_0(PE_wrapper321_U0_fifo_w_out_V_V_write_pass_0),
    .PE_wrapper322_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper322_U0_fifo_cout_drain_out_V_din_pass_0),
    .fifo_cout_drain_PE_14_4_V_full_n_pass_0(fifo_cout_drain_PE_14_4_V_full_n_pass_0),
    .PE_wrapper322_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper322_U0_fifo_cout_drain_out_V_write_pass_0),
    .cout_drain_IO_L1_out_wrapper401_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper401_U0_fifo_cout_drain_out_V_V_din_pass_0),
    .fifo_cout_drain_cout_drain_IO_L1_out_2_13_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_2_13_V_V_full_n_pass_0),
    .cout_drain_IO_L1_out_wrapper401_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper401_U0_fifo_cout_drain_out_V_V_write_pass_0),
    .cout_drain_IO_L1_out_wrapper434_U0_fifo_cout_drain_out_V_V_din_pass_0(cout_drain_IO_L1_out_wrapper434_U0_fifo_cout_drain_out_V_V_din_pass_0),
    .fifo_cout_drain_cout_drain_IO_L1_out_4_12_V_V_full_n_pass_0(fifo_cout_drain_cout_drain_IO_L1_out_4_12_V_V_full_n_pass_0),
    .cout_drain_IO_L1_out_wrapper434_U0_fifo_cout_drain_out_V_V_write_pass_0(cout_drain_IO_L1_out_wrapper434_U0_fifo_cout_drain_out_V_V_write_pass_0),
    .PE_wrapper298_U0_fifo_cout_drain_out_V_din_pass_0(PE_wrapper298_U0_fifo_cout_drain_out_V_din_pass_0),
    .fifo_cout_drain_PE_12_4_V_full_n_pass_0(fifo_cout_drain_PE_12_4_V_full_n_pass_0),
    .PE_wrapper298_U0_fifo_cout_drain_out_V_write_pass_0(PE_wrapper298_U0_fifo_cout_drain_out_V_write_pass_0),
    .ap_start(ap_start),
    .ap_done(ap_done),
    .ap_idle(ap_idle),
    .ap_ready(ap_ready),
    .ap_continue(ap_continue),
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n)
  );
endmodule


`timescale 1 ns / 1 ps


module CR_X2Y6_To_CR_X3Y7_routing (
input [31:0] PE_wrapper310_U0_fifo_cout_drain_out_V_din_pass_0,
output [31:0] PE_wrapper310_U0_fifo_cout_drain_out_V_din_pass_1,
output  fifo_cout_drain_PE_13_4_V_full_n_pass_0,
input  fifo_cout_drain_PE_13_4_V_full_n_pass_1,
input  PE_wrapper310_U0_fifo_cout_drain_out_V_write_pass_0,
output  PE_wrapper310_U0_fifo_cout_drain_out_V_write_pass_1,
input [31:0] PE_wrapper308_U0_fifo_cout_drain_out_V_din_pass_0,
output [31:0] PE_wrapper308_U0_fifo_cout_drain_out_V_din_pass_1,
output  fifo_cout_drain_PE_13_2_V_full_n_pass_0,
input  fifo_cout_drain_PE_13_2_V_full_n_pass_1,
input  PE_wrapper308_U0_fifo_cout_drain_out_V_write_pass_0,
output  PE_wrapper308_U0_fifo_cout_drain_out_V_write_pass_1,
input [255:0] PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0,
output [255:0] PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_1,
output  fifo_cin_PE_8_4_V_V_full_n_pass_0,
input  fifo_cin_PE_8_4_V_V_full_n_pass_1,
input  PE_wrapper238_U0_fifo_cin_out_V_V_write_pass_0,
output  PE_wrapper238_U0_fifo_cin_out_V_V_write_pass_1,
input [255:0] PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0,
output [255:0] PE_wrapper297_U0_fifo_w_out_V_V_din_pass_1,
output  fifo_w_PE_12_4_V_V_full_n_pass_0,
input  fifo_w_PE_12_4_V_V_full_n_pass_1,
input  PE_wrapper297_U0_fifo_w_out_V_V_write_pass_0,
output  PE_wrapper297_U0_fifo_w_out_V_V_write_pass_1,
input [255:0] PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0,
output [255:0] PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_1,
output  fifo_cin_PE_14_4_V_V_full_n_pass_0,
input  fifo_cin_PE_14_4_V_V_full_n_pass_1,
input  PE_wrapper310_U0_fifo_cin_out_V_V_write_pass_0,
output  PE_wrapper310_U0_fifo_cin_out_V_V_write_pass_1,
input [255:0] PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0,
output [255:0] PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_1,
output  fifo_cin_PE_14_1_V_V_full_n_pass_0,
input  fifo_cin_PE_14_1_V_V_full_n_pass_1,
input  PE_wrapper307_U0_fifo_cin_out_V_V_write_pass_0,
output  PE_wrapper307_U0_fifo_cin_out_V_V_write_pass_1,
input [255:0] PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0,
output [255:0] PE_wrapper250_U0_fifo_w_out_V_V_din_pass_1,
output  fifo_w_PE_8_5_V_V_full_n_pass_0,
input  fifo_w_PE_8_5_V_V_full_n_pass_1,
input  PE_wrapper250_U0_fifo_w_out_V_V_write_pass_0,
output  PE_wrapper250_U0_fifo_w_out_V_V_write_pass_1,
input [255:0] PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0,
output [255:0] PE_wrapper238_U0_fifo_w_out_V_V_din_pass_1,
output  fifo_w_PE_7_5_V_V_full_n_pass_0,
input  fifo_w_PE_7_5_V_V_full_n_pass_1,
input  PE_wrapper238_U0_fifo_w_out_V_V_write_pass_0,
output  PE_wrapper238_U0_fifo_w_out_V_V_write_pass_1,
output [31:0] PE_wrapper320_U0_fifo_cout_drain_out_V_din_pass_0,
input  fifo_cout_drain_PE_14_2_V_full_n_pass_0,
output  PE_wrapper320_U0_fifo_cout_drain_out_V_write_pass_0,
input [63:0] cout_drain_IO_L1_out_wrapper433_U0_fifo_cout_drain_out_V_V_din_pass_0,
output  fifo_cout_drain_cout_drain_IO_L1_out_4_13_V_V_full_n_pass_0,
input  cout_drain_IO_L1_out_wrapper433_U0_fifo_cout_drain_out_V_V_write_pass_0,
input [255:0] PE_wrapper309_U0_fifo_cin_out_V_V_din_pass_1,
output  fifo_cin_PE_14_3_V_V_full_n_pass_1,
input  PE_wrapper309_U0_fifo_cin_out_V_V_write_pass_1,
output [63:0] cout_drain_IO_L1_out_wrapper402_U0_fifo_cout_drain_out_V_V_din_pass_0,
input  fifo_cout_drain_cout_drain_IO_L1_out_2_12_V_V_full_n_pass_0,
output  cout_drain_IO_L1_out_wrapper402_U0_fifo_cout_drain_out_V_V_write_pass_0,
output [255:0] w_IO_L2_in149_U0_fifo_w_out_V_V_din_pass_0,
input  fifo_w_w_IO_L2_in_15_V_V_full_n_pass_0,
output  w_IO_L2_in149_U0_fifo_w_out_V_V_write_pass_0,
output [31:0] PE_wrapper286_U0_fifo_cout_drain_out_V_din_pass_0,
input  fifo_cout_drain_PE_11_4_V_full_n_pass_0,
output  PE_wrapper286_U0_fifo_cout_drain_out_V_write_pass_0,
input [255:0] PE_wrapper214_U0_fifo_cin_out_V_V_din_pass_1,
output  fifo_cin_PE_6_4_V_V_full_n_pass_1,
input  PE_wrapper214_U0_fifo_cin_out_V_V_write_pass_1,
output [63:0] cout_drain_IO_L1_out_wrapper432_U0_fifo_cout_drain_out_V_V_din_pass_0,
input  fifo_cout_drain_cout_drain_IO_L1_out_4_14_V_V_full_n_pass_0,
output  cout_drain_IO_L1_out_wrapper432_U0_fifo_cout_drain_out_V_V_write_pass_0,
output [255:0] PE_wrapper318_U0_fifo_w_out_V_V_din_pass_0,
input  fifo_w_PE_14_1_V_V_full_n_pass_0,
output  PE_wrapper318_U0_fifo_w_out_V_V_write_pass_0,
output [31:0] PE_wrapper226_U0_fifo_cout_drain_out_V_din_pass_0,
input  fifo_cout_drain_PE_6_4_V_full_n_pass_0,
output  PE_wrapper226_U0_fifo_cout_drain_out_V_write_pass_0,
output [255:0] PE_wrapper286_U0_fifo_cin_out_V_V_din_pass_0,
input  fifo_cin_PE_12_4_V_V_full_n_pass_0,
output  PE_wrapper286_U0_fifo_cin_out_V_V_write_pass_0,
input [255:0] w_IO_L2_in148_U0_fifo_w_out_V_V_din_pass_0,
output  fifo_w_w_IO_L2_in_14_V_V_full_n_pass_0,
input  w_IO_L2_in148_U0_fifo_w_out_V_V_write_pass_0,
output [255:0] PE_wrapper320_U0_fifo_cin_out_V_V_din_pass_0,
input  fifo_cin_PE_15_2_V_V_full_n_pass_0,
output  PE_wrapper320_U0_fifo_cin_out_V_V_write_pass_0,
input [63:0] cout_drain_IO_L1_out_wrapper418_U0_fifo_cout_drain_out_V_V_din_pass_1,
output  fifo_cout_drain_cout_drain_IO_L1_out_3_12_V_V_full_n_pass_1,
input  cout_drain_IO_L1_out_wrapper418_U0_fifo_cout_drain_out_V_V_write_pass_1,
input [255:0] PE_wrapper225_U0_fifo_w_out_V_V_din_pass_1,
output  fifo_w_PE_6_4_V_V_full_n_pass_1,
input  PE_wrapper225_U0_fifo_w_out_V_V_write_pass_1,
output [63:0] cout_drain_IO_L1_out_wrapper416_U0_fifo_cout_drain_out_V_V_din_pass_0,
input  fifo_cout_drain_cout_drain_IO_L1_out_3_14_V_V_full_n_pass_0,
output  cout_drain_IO_L1_out_wrapper416_U0_fifo_cout_drain_out_V_V_write_pass_0,
output [255:0] PE_wrapper330_U0_fifo_cin_out_V_V_din_pass_0,
input  fifo_cin_PE_16_0_V_V_full_n_pass_0,
output  PE_wrapper330_U0_fifo_cin_out_V_V_write_pass_0,
output [255:0] PE_wrapper330_U0_fifo_w_out_V_V_din_pass_0,
input  fifo_w_PE_15_1_V_V_full_n_pass_0,
output  PE_wrapper330_U0_fifo_w_out_V_V_write_pass_0,
input [255:0] PE_wrapper285_U0_fifo_w_out_V_V_din_pass_1,
output  fifo_w_PE_11_4_V_V_full_n_pass_1,
input  PE_wrapper285_U0_fifo_w_out_V_V_write_pass_1,
output [63:0] cout_drain_IO_L1_out_wrapper419_U0_fifo_cout_drain_out_V_V_din_pass_0,
input  fifo_cout_drain_cout_drain_IO_L1_out_3_11_V_V_full_n_pass_0,
output  cout_drain_IO_L1_out_wrapper419_U0_fifo_cout_drain_out_V_V_write_pass_0,
input [255:0] w_IO_L2_in_boundary_U0_fifo_w_local_out_V_V_din_pass_0,
output  fifo_w_PE_15_0_V_V_full_n_pass_0,
input  w_IO_L2_in_boundary_U0_fifo_w_local_out_V_V_write_pass_0,
input [255:0] PE_wrapper273_U0_fifo_w_out_V_V_din_pass_0,
output  fifo_w_PE_10_4_V_V_full_n_pass_0,
input  PE_wrapper273_U0_fifo_w_out_V_V_write_pass_0,
output [255:0] PE_wrapper286_U0_fifo_w_out_V_V_din_pass_0,
input  fifo_w_PE_11_5_V_V_full_n_pass_0,
output  PE_wrapper286_U0_fifo_w_out_V_V_write_pass_0,
input [63:0] cout_drain_IO_L1_out_boundary_wrapper383_U0_fifo_cout_drain_out_V_V_din_pass_0,
output  fifo_cout_drain_cout_drain_IO_L1_out_1_15_V_V_full_n_pass_0,
input  cout_drain_IO_L1_out_boundary_wrapper383_U0_fifo_cout_drain_out_V_V_write_pass_0,
output [31:0] PE_wrapper330_U0_fifo_cout_drain_out_V_din_pass_0,
input  fifo_cout_drain_PE_15_0_V_full_n_pass_0,
output  PE_wrapper330_U0_fifo_cout_drain_out_V_write_pass_0,
input [255:0] PE_wrapper306_U0_fifo_cin_out_V_V_din_pass_1,
output  fifo_cin_PE_14_0_V_V_full_n_pass_1,
input  PE_wrapper306_U0_fifo_cin_out_V_V_write_pass_1,
output [255:0] PE_wrapper321_U0_fifo_cin_out_V_V_din_pass_0,
input  fifo_cin_PE_15_3_V_V_full_n_pass_0,
output  PE_wrapper321_U0_fifo_cin_out_V_V_write_pass_0,
input [31:0] PE_wrapper285_U0_fifo_cout_drain_out_V_din_pass_1,
output  fifo_cout_drain_PE_11_3_V_full_n_pass_1,
input  PE_wrapper285_U0_fifo_cout_drain_out_V_write_pass_1,
input [255:0] PE_wrapper319_U0_fifo_w_out_V_V_din_pass_0,
output  fifo_w_PE_14_2_V_V_full_n_pass_0,
input  PE_wrapper319_U0_fifo_w_out_V_V_write_pass_0,
output [255:0] PE_wrapper226_U0_fifo_w_out_V_V_din_pass_0,
input  fifo_w_PE_6_5_V_V_full_n_pass_0,
output  PE_wrapper226_U0_fifo_w_out_V_V_write_pass_0,
input [255:0] PE_wrapper308_U0_fifo_cin_out_V_V_din_pass_0,
output  fifo_cin_PE_14_2_V_V_full_n_pass_0,
input  PE_wrapper308_U0_fifo_cin_out_V_V_write_pass_0,
output [63:0] cout_drain_IO_L1_out_wrapper384_U0_fifo_cout_drain_out_V_V_din_pass_0,
input  fifo_cout_drain_cout_drain_IO_L1_out_1_14_V_V_full_n_pass_0,
output  cout_drain_IO_L1_out_wrapper384_U0_fifo_cout_drain_out_V_V_write_pass_0,
input [31:0] PE_wrapper319_U0_fifo_cout_drain_out_V_din_pass_0,
output  fifo_cout_drain_PE_14_1_V_full_n_pass_0,
input  PE_wrapper319_U0_fifo_cout_drain_out_V_write_pass_0,
input [31:0] PE_wrapper334_U0_fifo_cout_drain_out_V_din_pass_0,
output  fifo_cout_drain_PE_15_4_V_full_n_pass_0,
input  PE_wrapper334_U0_fifo_cout_drain_out_V_write_pass_0,
input [63:0] cout_drain_IO_L1_out_boundary_wrapper415_U0_fifo_cout_drain_out_V_V_din_pass_0,
output  fifo_cout_drain_cout_drain_IO_L1_out_3_15_V_V_full_n_pass_0,
input  cout_drain_IO_L1_out_boundary_wrapper415_U0_fifo_cout_drain_out_V_V_write_pass_0,
output [255:0] PE_wrapper274_U0_fifo_w_out_V_V_din_pass_0,
input  fifo_w_PE_10_5_V_V_full_n_pass_0,
output  PE_wrapper274_U0_fifo_w_out_V_V_write_pass_0,
input [255:0] PE_wrapper262_U0_fifo_cin_out_V_V_din_pass_1,
output  fifo_cin_PE_10_4_V_V_full_n_pass_1,
input  PE_wrapper262_U0_fifo_cin_out_V_V_write_pass_1,
output [255:0] PE_wrapper226_U0_fifo_cin_out_V_V_din_pass_0,
input  fifo_cin_PE_7_4_V_V_full_n_pass_0,
output  PE_wrapper226_U0_fifo_cin_out_V_V_write_pass_0,
output [31:0] PE_wrapper318_U0_fifo_cout_drain_out_V_din_pass_0,
input  fifo_cout_drain_PE_14_0_V_full_n_pass_0,
output  PE_wrapper318_U0_fifo_cout_drain_out_V_write_pass_0,
output [31:0] PE_wrapper274_U0_fifo_cout_drain_out_V_din_pass_0,
input  fifo_cout_drain_PE_10_4_V_full_n_pass_0,
output  PE_wrapper274_U0_fifo_cout_drain_out_V_write_pass_0,
input [31:0] PE_wrapper296_U0_fifo_cout_drain_out_V_din_pass_1,
output  fifo_cout_drain_PE_12_2_V_full_n_pass_1,
input  PE_wrapper296_U0_fifo_cout_drain_out_V_write_pass_1,
output [255:0] PE_wrapper321_U0_fifo_w_out_V_V_din_pass_0,
input  fifo_w_PE_14_4_V_V_full_n_pass_0,
output  PE_wrapper321_U0_fifo_w_out_V_V_write_pass_0,
input [31:0] PE_wrapper322_U0_fifo_cout_drain_out_V_din_pass_0,
output  fifo_cout_drain_PE_14_4_V_full_n_pass_0,
input  PE_wrapper322_U0_fifo_cout_drain_out_V_write_pass_0,
input [63:0] cout_drain_IO_L1_out_wrapper401_U0_fifo_cout_drain_out_V_V_din_pass_0,
output  fifo_cout_drain_cout_drain_IO_L1_out_2_13_V_V_full_n_pass_0,
input  cout_drain_IO_L1_out_wrapper401_U0_fifo_cout_drain_out_V_V_write_pass_0,
output [63:0] cout_drain_IO_L1_out_wrapper434_U0_fifo_cout_drain_out_V_V_din_pass_0,
input  fifo_cout_drain_cout_drain_IO_L1_out_4_12_V_V_full_n_pass_0,
output  cout_drain_IO_L1_out_wrapper434_U0_fifo_cout_drain_out_V_V_write_pass_0,
input [31:0] PE_wrapper298_U0_fifo_cout_drain_out_V_din_pass_0,
output  fifo_cout_drain_PE_12_4_V_full_n_pass_0,
input  PE_wrapper298_U0_fifo_cout_drain_out_V_write_pass_0,
input ap_start,
output ap_done,
output ap_idle,
output ap_ready,
input ap_continue,
input ap_clk,
input ap_rst_n
);
  wire [31:0] PE_wrapper310_U0_fifo_cout_drain_out_V_din_q0;
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cout_drain_out_V_din_q0_0_lut ( .O(PE_wrapper310_U0_fifo_cout_drain_out_V_din_q0[0]), .I0(PE_wrapper310_U0_fifo_cout_drain_out_V_din_pass_0[0]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cout_drain_out_V_din_q0_1_lut ( .O(PE_wrapper310_U0_fifo_cout_drain_out_V_din_q0[1]), .I0(PE_wrapper310_U0_fifo_cout_drain_out_V_din_pass_0[1]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cout_drain_out_V_din_q0_2_lut ( .O(PE_wrapper310_U0_fifo_cout_drain_out_V_din_q0[2]), .I0(PE_wrapper310_U0_fifo_cout_drain_out_V_din_pass_0[2]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cout_drain_out_V_din_q0_3_lut ( .O(PE_wrapper310_U0_fifo_cout_drain_out_V_din_q0[3]), .I0(PE_wrapper310_U0_fifo_cout_drain_out_V_din_pass_0[3]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cout_drain_out_V_din_q0_4_lut ( .O(PE_wrapper310_U0_fifo_cout_drain_out_V_din_q0[4]), .I0(PE_wrapper310_U0_fifo_cout_drain_out_V_din_pass_0[4]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cout_drain_out_V_din_q0_5_lut ( .O(PE_wrapper310_U0_fifo_cout_drain_out_V_din_q0[5]), .I0(PE_wrapper310_U0_fifo_cout_drain_out_V_din_pass_0[5]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cout_drain_out_V_din_q0_6_lut ( .O(PE_wrapper310_U0_fifo_cout_drain_out_V_din_q0[6]), .I0(PE_wrapper310_U0_fifo_cout_drain_out_V_din_pass_0[6]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cout_drain_out_V_din_q0_7_lut ( .O(PE_wrapper310_U0_fifo_cout_drain_out_V_din_q0[7]), .I0(PE_wrapper310_U0_fifo_cout_drain_out_V_din_pass_0[7]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cout_drain_out_V_din_q0_8_lut ( .O(PE_wrapper310_U0_fifo_cout_drain_out_V_din_q0[8]), .I0(PE_wrapper310_U0_fifo_cout_drain_out_V_din_pass_0[8]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cout_drain_out_V_din_q0_9_lut ( .O(PE_wrapper310_U0_fifo_cout_drain_out_V_din_q0[9]), .I0(PE_wrapper310_U0_fifo_cout_drain_out_V_din_pass_0[9]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cout_drain_out_V_din_q0_10_lut ( .O(PE_wrapper310_U0_fifo_cout_drain_out_V_din_q0[10]), .I0(PE_wrapper310_U0_fifo_cout_drain_out_V_din_pass_0[10]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cout_drain_out_V_din_q0_11_lut ( .O(PE_wrapper310_U0_fifo_cout_drain_out_V_din_q0[11]), .I0(PE_wrapper310_U0_fifo_cout_drain_out_V_din_pass_0[11]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cout_drain_out_V_din_q0_12_lut ( .O(PE_wrapper310_U0_fifo_cout_drain_out_V_din_q0[12]), .I0(PE_wrapper310_U0_fifo_cout_drain_out_V_din_pass_0[12]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cout_drain_out_V_din_q0_13_lut ( .O(PE_wrapper310_U0_fifo_cout_drain_out_V_din_q0[13]), .I0(PE_wrapper310_U0_fifo_cout_drain_out_V_din_pass_0[13]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cout_drain_out_V_din_q0_14_lut ( .O(PE_wrapper310_U0_fifo_cout_drain_out_V_din_q0[14]), .I0(PE_wrapper310_U0_fifo_cout_drain_out_V_din_pass_0[14]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cout_drain_out_V_din_q0_15_lut ( .O(PE_wrapper310_U0_fifo_cout_drain_out_V_din_q0[15]), .I0(PE_wrapper310_U0_fifo_cout_drain_out_V_din_pass_0[15]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cout_drain_out_V_din_q0_16_lut ( .O(PE_wrapper310_U0_fifo_cout_drain_out_V_din_q0[16]), .I0(PE_wrapper310_U0_fifo_cout_drain_out_V_din_pass_0[16]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cout_drain_out_V_din_q0_17_lut ( .O(PE_wrapper310_U0_fifo_cout_drain_out_V_din_q0[17]), .I0(PE_wrapper310_U0_fifo_cout_drain_out_V_din_pass_0[17]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cout_drain_out_V_din_q0_18_lut ( .O(PE_wrapper310_U0_fifo_cout_drain_out_V_din_q0[18]), .I0(PE_wrapper310_U0_fifo_cout_drain_out_V_din_pass_0[18]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cout_drain_out_V_din_q0_19_lut ( .O(PE_wrapper310_U0_fifo_cout_drain_out_V_din_q0[19]), .I0(PE_wrapper310_U0_fifo_cout_drain_out_V_din_pass_0[19]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cout_drain_out_V_din_q0_20_lut ( .O(PE_wrapper310_U0_fifo_cout_drain_out_V_din_q0[20]), .I0(PE_wrapper310_U0_fifo_cout_drain_out_V_din_pass_0[20]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cout_drain_out_V_din_q0_21_lut ( .O(PE_wrapper310_U0_fifo_cout_drain_out_V_din_q0[21]), .I0(PE_wrapper310_U0_fifo_cout_drain_out_V_din_pass_0[21]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cout_drain_out_V_din_q0_22_lut ( .O(PE_wrapper310_U0_fifo_cout_drain_out_V_din_q0[22]), .I0(PE_wrapper310_U0_fifo_cout_drain_out_V_din_pass_0[22]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cout_drain_out_V_din_q0_23_lut ( .O(PE_wrapper310_U0_fifo_cout_drain_out_V_din_q0[23]), .I0(PE_wrapper310_U0_fifo_cout_drain_out_V_din_pass_0[23]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cout_drain_out_V_din_q0_24_lut ( .O(PE_wrapper310_U0_fifo_cout_drain_out_V_din_q0[24]), .I0(PE_wrapper310_U0_fifo_cout_drain_out_V_din_pass_0[24]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cout_drain_out_V_din_q0_25_lut ( .O(PE_wrapper310_U0_fifo_cout_drain_out_V_din_q0[25]), .I0(PE_wrapper310_U0_fifo_cout_drain_out_V_din_pass_0[25]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cout_drain_out_V_din_q0_26_lut ( .O(PE_wrapper310_U0_fifo_cout_drain_out_V_din_q0[26]), .I0(PE_wrapper310_U0_fifo_cout_drain_out_V_din_pass_0[26]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cout_drain_out_V_din_q0_27_lut ( .O(PE_wrapper310_U0_fifo_cout_drain_out_V_din_q0[27]), .I0(PE_wrapper310_U0_fifo_cout_drain_out_V_din_pass_0[27]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cout_drain_out_V_din_q0_28_lut ( .O(PE_wrapper310_U0_fifo_cout_drain_out_V_din_q0[28]), .I0(PE_wrapper310_U0_fifo_cout_drain_out_V_din_pass_0[28]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cout_drain_out_V_din_q0_29_lut ( .O(PE_wrapper310_U0_fifo_cout_drain_out_V_din_q0[29]), .I0(PE_wrapper310_U0_fifo_cout_drain_out_V_din_pass_0[29]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cout_drain_out_V_din_q0_30_lut ( .O(PE_wrapper310_U0_fifo_cout_drain_out_V_din_q0[30]), .I0(PE_wrapper310_U0_fifo_cout_drain_out_V_din_pass_0[30]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cout_drain_out_V_din_q0_31_lut ( .O(PE_wrapper310_U0_fifo_cout_drain_out_V_din_q0[31]), .I0(PE_wrapper310_U0_fifo_cout_drain_out_V_din_pass_0[31]) );
  assign PE_wrapper310_U0_fifo_cout_drain_out_V_din_pass_1 = PE_wrapper310_U0_fifo_cout_drain_out_V_din_q0;
  wire  fifo_cout_drain_PE_13_4_V_full_n_q0;
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) fifo_cout_drain_PE_13_4_V_full_n_q0_lut ( .O(fifo_cout_drain_PE_13_4_V_full_n_q0), .I0(fifo_cout_drain_PE_13_4_V_full_n_pass_1) );
  assign fifo_cout_drain_PE_13_4_V_full_n_pass_0 = fifo_cout_drain_PE_13_4_V_full_n_q0;
  wire  PE_wrapper310_U0_fifo_cout_drain_out_V_write_q0;
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cout_drain_out_V_write_q0_lut ( .O(PE_wrapper310_U0_fifo_cout_drain_out_V_write_q0), .I0(PE_wrapper310_U0_fifo_cout_drain_out_V_write_pass_0) );
  assign PE_wrapper310_U0_fifo_cout_drain_out_V_write_pass_1 = PE_wrapper310_U0_fifo_cout_drain_out_V_write_q0;
  wire [31:0] PE_wrapper308_U0_fifo_cout_drain_out_V_din_q0;
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper308_U0_fifo_cout_drain_out_V_din_q0_0_lut ( .O(PE_wrapper308_U0_fifo_cout_drain_out_V_din_q0[0]), .I0(PE_wrapper308_U0_fifo_cout_drain_out_V_din_pass_0[0]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper308_U0_fifo_cout_drain_out_V_din_q0_1_lut ( .O(PE_wrapper308_U0_fifo_cout_drain_out_V_din_q0[1]), .I0(PE_wrapper308_U0_fifo_cout_drain_out_V_din_pass_0[1]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper308_U0_fifo_cout_drain_out_V_din_q0_2_lut ( .O(PE_wrapper308_U0_fifo_cout_drain_out_V_din_q0[2]), .I0(PE_wrapper308_U0_fifo_cout_drain_out_V_din_pass_0[2]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper308_U0_fifo_cout_drain_out_V_din_q0_3_lut ( .O(PE_wrapper308_U0_fifo_cout_drain_out_V_din_q0[3]), .I0(PE_wrapper308_U0_fifo_cout_drain_out_V_din_pass_0[3]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper308_U0_fifo_cout_drain_out_V_din_q0_4_lut ( .O(PE_wrapper308_U0_fifo_cout_drain_out_V_din_q0[4]), .I0(PE_wrapper308_U0_fifo_cout_drain_out_V_din_pass_0[4]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper308_U0_fifo_cout_drain_out_V_din_q0_5_lut ( .O(PE_wrapper308_U0_fifo_cout_drain_out_V_din_q0[5]), .I0(PE_wrapper308_U0_fifo_cout_drain_out_V_din_pass_0[5]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper308_U0_fifo_cout_drain_out_V_din_q0_6_lut ( .O(PE_wrapper308_U0_fifo_cout_drain_out_V_din_q0[6]), .I0(PE_wrapper308_U0_fifo_cout_drain_out_V_din_pass_0[6]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper308_U0_fifo_cout_drain_out_V_din_q0_7_lut ( .O(PE_wrapper308_U0_fifo_cout_drain_out_V_din_q0[7]), .I0(PE_wrapper308_U0_fifo_cout_drain_out_V_din_pass_0[7]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper308_U0_fifo_cout_drain_out_V_din_q0_8_lut ( .O(PE_wrapper308_U0_fifo_cout_drain_out_V_din_q0[8]), .I0(PE_wrapper308_U0_fifo_cout_drain_out_V_din_pass_0[8]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper308_U0_fifo_cout_drain_out_V_din_q0_9_lut ( .O(PE_wrapper308_U0_fifo_cout_drain_out_V_din_q0[9]), .I0(PE_wrapper308_U0_fifo_cout_drain_out_V_din_pass_0[9]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper308_U0_fifo_cout_drain_out_V_din_q0_10_lut ( .O(PE_wrapper308_U0_fifo_cout_drain_out_V_din_q0[10]), .I0(PE_wrapper308_U0_fifo_cout_drain_out_V_din_pass_0[10]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper308_U0_fifo_cout_drain_out_V_din_q0_11_lut ( .O(PE_wrapper308_U0_fifo_cout_drain_out_V_din_q0[11]), .I0(PE_wrapper308_U0_fifo_cout_drain_out_V_din_pass_0[11]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper308_U0_fifo_cout_drain_out_V_din_q0_12_lut ( .O(PE_wrapper308_U0_fifo_cout_drain_out_V_din_q0[12]), .I0(PE_wrapper308_U0_fifo_cout_drain_out_V_din_pass_0[12]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper308_U0_fifo_cout_drain_out_V_din_q0_13_lut ( .O(PE_wrapper308_U0_fifo_cout_drain_out_V_din_q0[13]), .I0(PE_wrapper308_U0_fifo_cout_drain_out_V_din_pass_0[13]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper308_U0_fifo_cout_drain_out_V_din_q0_14_lut ( .O(PE_wrapper308_U0_fifo_cout_drain_out_V_din_q0[14]), .I0(PE_wrapper308_U0_fifo_cout_drain_out_V_din_pass_0[14]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper308_U0_fifo_cout_drain_out_V_din_q0_15_lut ( .O(PE_wrapper308_U0_fifo_cout_drain_out_V_din_q0[15]), .I0(PE_wrapper308_U0_fifo_cout_drain_out_V_din_pass_0[15]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper308_U0_fifo_cout_drain_out_V_din_q0_16_lut ( .O(PE_wrapper308_U0_fifo_cout_drain_out_V_din_q0[16]), .I0(PE_wrapper308_U0_fifo_cout_drain_out_V_din_pass_0[16]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper308_U0_fifo_cout_drain_out_V_din_q0_17_lut ( .O(PE_wrapper308_U0_fifo_cout_drain_out_V_din_q0[17]), .I0(PE_wrapper308_U0_fifo_cout_drain_out_V_din_pass_0[17]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper308_U0_fifo_cout_drain_out_V_din_q0_18_lut ( .O(PE_wrapper308_U0_fifo_cout_drain_out_V_din_q0[18]), .I0(PE_wrapper308_U0_fifo_cout_drain_out_V_din_pass_0[18]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper308_U0_fifo_cout_drain_out_V_din_q0_19_lut ( .O(PE_wrapper308_U0_fifo_cout_drain_out_V_din_q0[19]), .I0(PE_wrapper308_U0_fifo_cout_drain_out_V_din_pass_0[19]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper308_U0_fifo_cout_drain_out_V_din_q0_20_lut ( .O(PE_wrapper308_U0_fifo_cout_drain_out_V_din_q0[20]), .I0(PE_wrapper308_U0_fifo_cout_drain_out_V_din_pass_0[20]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper308_U0_fifo_cout_drain_out_V_din_q0_21_lut ( .O(PE_wrapper308_U0_fifo_cout_drain_out_V_din_q0[21]), .I0(PE_wrapper308_U0_fifo_cout_drain_out_V_din_pass_0[21]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper308_U0_fifo_cout_drain_out_V_din_q0_22_lut ( .O(PE_wrapper308_U0_fifo_cout_drain_out_V_din_q0[22]), .I0(PE_wrapper308_U0_fifo_cout_drain_out_V_din_pass_0[22]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper308_U0_fifo_cout_drain_out_V_din_q0_23_lut ( .O(PE_wrapper308_U0_fifo_cout_drain_out_V_din_q0[23]), .I0(PE_wrapper308_U0_fifo_cout_drain_out_V_din_pass_0[23]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper308_U0_fifo_cout_drain_out_V_din_q0_24_lut ( .O(PE_wrapper308_U0_fifo_cout_drain_out_V_din_q0[24]), .I0(PE_wrapper308_U0_fifo_cout_drain_out_V_din_pass_0[24]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper308_U0_fifo_cout_drain_out_V_din_q0_25_lut ( .O(PE_wrapper308_U0_fifo_cout_drain_out_V_din_q0[25]), .I0(PE_wrapper308_U0_fifo_cout_drain_out_V_din_pass_0[25]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper308_U0_fifo_cout_drain_out_V_din_q0_26_lut ( .O(PE_wrapper308_U0_fifo_cout_drain_out_V_din_q0[26]), .I0(PE_wrapper308_U0_fifo_cout_drain_out_V_din_pass_0[26]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper308_U0_fifo_cout_drain_out_V_din_q0_27_lut ( .O(PE_wrapper308_U0_fifo_cout_drain_out_V_din_q0[27]), .I0(PE_wrapper308_U0_fifo_cout_drain_out_V_din_pass_0[27]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper308_U0_fifo_cout_drain_out_V_din_q0_28_lut ( .O(PE_wrapper308_U0_fifo_cout_drain_out_V_din_q0[28]), .I0(PE_wrapper308_U0_fifo_cout_drain_out_V_din_pass_0[28]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper308_U0_fifo_cout_drain_out_V_din_q0_29_lut ( .O(PE_wrapper308_U0_fifo_cout_drain_out_V_din_q0[29]), .I0(PE_wrapper308_U0_fifo_cout_drain_out_V_din_pass_0[29]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper308_U0_fifo_cout_drain_out_V_din_q0_30_lut ( .O(PE_wrapper308_U0_fifo_cout_drain_out_V_din_q0[30]), .I0(PE_wrapper308_U0_fifo_cout_drain_out_V_din_pass_0[30]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper308_U0_fifo_cout_drain_out_V_din_q0_31_lut ( .O(PE_wrapper308_U0_fifo_cout_drain_out_V_din_q0[31]), .I0(PE_wrapper308_U0_fifo_cout_drain_out_V_din_pass_0[31]) );
  assign PE_wrapper308_U0_fifo_cout_drain_out_V_din_pass_1 = PE_wrapper308_U0_fifo_cout_drain_out_V_din_q0;
  wire  fifo_cout_drain_PE_13_2_V_full_n_q0;
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) fifo_cout_drain_PE_13_2_V_full_n_q0_lut ( .O(fifo_cout_drain_PE_13_2_V_full_n_q0), .I0(fifo_cout_drain_PE_13_2_V_full_n_pass_1) );
  assign fifo_cout_drain_PE_13_2_V_full_n_pass_0 = fifo_cout_drain_PE_13_2_V_full_n_q0;
  wire  PE_wrapper308_U0_fifo_cout_drain_out_V_write_q0;
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper308_U0_fifo_cout_drain_out_V_write_q0_lut ( .O(PE_wrapper308_U0_fifo_cout_drain_out_V_write_q0), .I0(PE_wrapper308_U0_fifo_cout_drain_out_V_write_pass_0) );
  assign PE_wrapper308_U0_fifo_cout_drain_out_V_write_pass_1 = PE_wrapper308_U0_fifo_cout_drain_out_V_write_q0;
  wire [255:0] PE_wrapper238_U0_fifo_cin_out_V_V_din_q0;
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_0_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[0]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[0]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_1_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[1]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[1]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_2_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[2]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[2]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_3_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[3]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[3]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_4_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[4]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[4]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_5_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[5]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[5]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_6_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[6]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[6]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_7_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[7]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[7]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_8_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[8]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[8]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_9_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[9]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[9]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_10_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[10]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[10]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_11_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[11]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[11]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_12_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[12]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[12]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_13_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[13]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[13]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_14_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[14]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[14]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_15_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[15]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[15]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_16_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[16]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[16]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_17_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[17]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[17]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_18_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[18]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[18]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_19_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[19]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[19]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_20_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[20]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[20]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_21_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[21]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[21]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_22_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[22]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[22]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_23_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[23]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[23]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_24_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[24]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[24]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_25_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[25]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[25]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_26_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[26]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[26]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_27_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[27]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[27]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_28_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[28]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[28]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_29_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[29]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[29]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_30_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[30]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[30]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_31_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[31]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[31]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_32_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[32]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[32]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_33_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[33]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[33]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_34_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[34]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[34]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_35_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[35]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[35]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_36_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[36]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[36]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_37_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[37]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[37]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_38_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[38]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[38]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_39_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[39]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[39]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_40_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[40]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[40]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_41_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[41]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[41]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_42_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[42]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[42]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_43_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[43]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[43]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_44_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[44]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[44]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_45_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[45]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[45]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_46_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[46]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[46]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_47_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[47]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[47]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_48_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[48]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[48]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_49_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[49]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[49]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_50_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[50]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[50]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_51_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[51]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[51]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_52_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[52]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[52]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_53_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[53]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[53]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_54_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[54]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[54]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_55_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[55]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[55]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_56_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[56]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[56]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_57_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[57]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[57]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_58_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[58]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[58]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_59_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[59]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[59]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_60_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[60]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[60]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_61_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[61]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[61]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_62_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[62]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[62]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_63_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[63]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[63]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_64_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[64]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[64]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_65_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[65]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[65]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_66_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[66]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[66]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_67_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[67]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[67]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_68_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[68]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[68]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_69_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[69]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[69]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_70_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[70]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[70]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_71_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[71]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[71]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_72_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[72]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[72]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_73_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[73]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[73]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_74_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[74]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[74]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_75_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[75]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[75]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_76_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[76]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[76]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_77_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[77]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[77]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_78_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[78]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[78]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_79_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[79]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[79]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_80_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[80]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[80]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_81_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[81]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[81]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_82_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[82]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[82]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_83_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[83]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[83]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_84_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[84]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[84]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_85_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[85]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[85]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_86_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[86]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[86]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_87_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[87]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[87]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_88_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[88]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[88]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_89_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[89]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[89]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_90_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[90]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[90]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_91_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[91]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[91]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_92_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[92]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[92]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_93_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[93]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[93]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_94_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[94]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[94]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_95_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[95]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[95]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_96_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[96]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[96]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_97_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[97]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[97]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_98_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[98]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[98]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_99_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[99]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[99]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_100_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[100]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[100]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_101_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[101]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[101]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_102_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[102]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[102]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_103_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[103]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[103]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_104_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[104]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[104]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_105_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[105]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[105]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_106_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[106]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[106]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_107_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[107]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[107]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_108_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[108]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[108]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_109_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[109]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[109]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_110_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[110]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[110]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_111_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[111]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[111]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_112_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[112]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[112]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_113_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[113]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[113]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_114_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[114]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[114]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_115_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[115]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[115]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_116_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[116]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[116]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_117_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[117]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[117]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_118_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[118]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[118]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_119_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[119]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[119]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_120_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[120]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[120]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_121_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[121]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[121]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_122_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[122]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[122]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_123_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[123]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[123]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_124_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[124]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[124]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_125_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[125]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[125]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_126_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[126]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[126]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_127_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[127]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[127]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_128_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[128]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[128]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_129_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[129]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[129]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_130_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[130]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[130]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_131_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[131]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[131]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_132_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[132]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[132]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_133_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[133]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[133]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_134_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[134]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[134]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_135_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[135]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[135]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_136_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[136]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[136]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_137_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[137]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[137]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_138_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[138]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[138]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_139_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[139]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[139]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_140_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[140]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[140]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_141_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[141]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[141]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_142_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[142]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[142]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_143_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[143]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[143]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_144_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[144]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[144]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_145_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[145]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[145]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_146_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[146]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[146]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_147_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[147]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[147]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_148_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[148]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[148]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_149_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[149]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[149]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_150_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[150]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[150]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_151_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[151]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[151]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_152_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[152]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[152]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_153_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[153]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[153]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_154_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[154]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[154]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_155_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[155]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[155]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_156_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[156]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[156]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_157_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[157]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[157]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_158_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[158]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[158]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_159_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[159]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[159]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_160_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[160]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[160]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_161_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[161]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[161]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_162_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[162]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[162]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_163_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[163]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[163]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_164_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[164]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[164]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_165_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[165]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[165]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_166_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[166]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[166]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_167_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[167]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[167]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_168_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[168]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[168]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_169_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[169]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[169]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_170_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[170]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[170]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_171_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[171]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[171]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_172_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[172]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[172]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_173_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[173]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[173]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_174_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[174]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[174]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_175_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[175]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[175]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_176_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[176]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[176]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_177_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[177]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[177]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_178_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[178]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[178]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_179_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[179]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[179]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_180_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[180]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[180]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_181_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[181]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[181]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_182_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[182]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[182]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_183_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[183]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[183]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_184_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[184]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[184]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_185_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[185]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[185]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_186_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[186]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[186]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_187_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[187]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[187]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_188_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[188]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[188]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_189_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[189]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[189]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_190_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[190]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[190]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_191_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[191]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[191]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_192_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[192]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[192]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_193_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[193]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[193]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_194_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[194]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[194]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_195_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[195]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[195]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_196_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[196]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[196]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_197_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[197]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[197]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_198_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[198]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[198]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_199_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[199]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[199]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_200_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[200]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[200]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_201_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[201]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[201]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_202_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[202]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[202]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_203_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[203]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[203]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_204_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[204]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[204]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_205_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[205]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[205]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_206_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[206]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[206]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_207_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[207]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[207]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_208_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[208]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[208]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_209_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[209]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[209]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_210_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[210]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[210]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_211_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[211]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[211]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_212_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[212]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[212]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_213_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[213]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[213]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_214_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[214]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[214]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_215_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[215]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[215]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_216_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[216]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[216]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_217_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[217]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[217]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_218_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[218]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[218]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_219_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[219]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[219]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_220_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[220]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[220]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_221_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[221]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[221]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_222_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[222]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[222]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_223_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[223]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[223]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_224_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[224]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[224]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_225_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[225]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[225]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_226_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[226]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[226]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_227_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[227]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[227]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_228_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[228]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[228]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_229_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[229]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[229]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_230_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[230]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[230]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_231_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[231]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[231]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_232_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[232]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[232]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_233_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[233]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[233]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_234_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[234]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[234]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_235_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[235]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[235]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_236_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[236]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[236]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_237_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[237]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[237]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_238_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[238]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[238]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_239_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[239]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[239]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_240_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[240]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[240]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_241_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[241]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[241]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_242_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[242]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[242]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_243_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[243]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[243]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_244_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[244]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[244]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_245_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[245]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[245]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_246_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[246]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[246]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_247_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[247]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[247]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_248_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[248]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[248]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_249_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[249]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[249]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_250_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[250]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[250]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_251_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[251]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[251]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_252_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[252]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[252]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_253_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[253]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[253]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_254_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[254]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[254]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_din_q0_255_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_din_q0[255]), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_0[255]) );
  assign PE_wrapper238_U0_fifo_cin_out_V_V_din_pass_1 = PE_wrapper238_U0_fifo_cin_out_V_V_din_q0;
  wire  fifo_cin_PE_8_4_V_V_full_n_q0;
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) fifo_cin_PE_8_4_V_V_full_n_q0_lut ( .O(fifo_cin_PE_8_4_V_V_full_n_q0), .I0(fifo_cin_PE_8_4_V_V_full_n_pass_1) );
  assign fifo_cin_PE_8_4_V_V_full_n_pass_0 = fifo_cin_PE_8_4_V_V_full_n_q0;
  wire  PE_wrapper238_U0_fifo_cin_out_V_V_write_q0;
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_cin_out_V_V_write_q0_lut ( .O(PE_wrapper238_U0_fifo_cin_out_V_V_write_q0), .I0(PE_wrapper238_U0_fifo_cin_out_V_V_write_pass_0) );
  assign PE_wrapper238_U0_fifo_cin_out_V_V_write_pass_1 = PE_wrapper238_U0_fifo_cin_out_V_V_write_q0;
  wire [255:0] PE_wrapper297_U0_fifo_w_out_V_V_din_q0;
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_0_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[0]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[0]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_1_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[1]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[1]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_2_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[2]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[2]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_3_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[3]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[3]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_4_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[4]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[4]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_5_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[5]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[5]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_6_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[6]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[6]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_7_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[7]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[7]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_8_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[8]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[8]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_9_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[9]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[9]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_10_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[10]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[10]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_11_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[11]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[11]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_12_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[12]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[12]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_13_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[13]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[13]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_14_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[14]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[14]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_15_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[15]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[15]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_16_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[16]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[16]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_17_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[17]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[17]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_18_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[18]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[18]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_19_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[19]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[19]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_20_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[20]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[20]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_21_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[21]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[21]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_22_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[22]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[22]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_23_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[23]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[23]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_24_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[24]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[24]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_25_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[25]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[25]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_26_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[26]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[26]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_27_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[27]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[27]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_28_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[28]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[28]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_29_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[29]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[29]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_30_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[30]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[30]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_31_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[31]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[31]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_32_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[32]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[32]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_33_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[33]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[33]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_34_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[34]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[34]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_35_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[35]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[35]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_36_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[36]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[36]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_37_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[37]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[37]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_38_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[38]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[38]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_39_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[39]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[39]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_40_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[40]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[40]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_41_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[41]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[41]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_42_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[42]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[42]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_43_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[43]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[43]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_44_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[44]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[44]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_45_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[45]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[45]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_46_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[46]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[46]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_47_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[47]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[47]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_48_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[48]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[48]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_49_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[49]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[49]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_50_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[50]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[50]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_51_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[51]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[51]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_52_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[52]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[52]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_53_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[53]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[53]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_54_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[54]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[54]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_55_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[55]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[55]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_56_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[56]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[56]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_57_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[57]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[57]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_58_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[58]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[58]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_59_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[59]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[59]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_60_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[60]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[60]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_61_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[61]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[61]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_62_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[62]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[62]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_63_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[63]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[63]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_64_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[64]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[64]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_65_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[65]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[65]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_66_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[66]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[66]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_67_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[67]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[67]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_68_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[68]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[68]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_69_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[69]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[69]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_70_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[70]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[70]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_71_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[71]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[71]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_72_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[72]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[72]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_73_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[73]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[73]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_74_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[74]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[74]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_75_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[75]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[75]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_76_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[76]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[76]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_77_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[77]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[77]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_78_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[78]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[78]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_79_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[79]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[79]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_80_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[80]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[80]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_81_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[81]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[81]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_82_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[82]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[82]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_83_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[83]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[83]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_84_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[84]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[84]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_85_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[85]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[85]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_86_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[86]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[86]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_87_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[87]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[87]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_88_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[88]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[88]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_89_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[89]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[89]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_90_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[90]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[90]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_91_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[91]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[91]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_92_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[92]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[92]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_93_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[93]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[93]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_94_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[94]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[94]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_95_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[95]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[95]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_96_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[96]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[96]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_97_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[97]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[97]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_98_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[98]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[98]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_99_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[99]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[99]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_100_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[100]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[100]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_101_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[101]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[101]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_102_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[102]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[102]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_103_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[103]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[103]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_104_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[104]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[104]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_105_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[105]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[105]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_106_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[106]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[106]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_107_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[107]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[107]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_108_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[108]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[108]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_109_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[109]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[109]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_110_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[110]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[110]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_111_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[111]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[111]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_112_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[112]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[112]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_113_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[113]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[113]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_114_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[114]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[114]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_115_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[115]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[115]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_116_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[116]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[116]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_117_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[117]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[117]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_118_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[118]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[118]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_119_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[119]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[119]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_120_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[120]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[120]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_121_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[121]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[121]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_122_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[122]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[122]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_123_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[123]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[123]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_124_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[124]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[124]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_125_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[125]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[125]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_126_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[126]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[126]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_127_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[127]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[127]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_128_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[128]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[128]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_129_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[129]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[129]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_130_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[130]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[130]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_131_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[131]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[131]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_132_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[132]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[132]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_133_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[133]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[133]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_134_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[134]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[134]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_135_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[135]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[135]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_136_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[136]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[136]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_137_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[137]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[137]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_138_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[138]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[138]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_139_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[139]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[139]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_140_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[140]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[140]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_141_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[141]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[141]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_142_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[142]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[142]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_143_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[143]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[143]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_144_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[144]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[144]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_145_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[145]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[145]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_146_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[146]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[146]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_147_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[147]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[147]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_148_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[148]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[148]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_149_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[149]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[149]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_150_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[150]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[150]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_151_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[151]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[151]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_152_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[152]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[152]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_153_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[153]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[153]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_154_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[154]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[154]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_155_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[155]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[155]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_156_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[156]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[156]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_157_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[157]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[157]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_158_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[158]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[158]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_159_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[159]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[159]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_160_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[160]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[160]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_161_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[161]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[161]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_162_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[162]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[162]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_163_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[163]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[163]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_164_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[164]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[164]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_165_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[165]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[165]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_166_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[166]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[166]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_167_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[167]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[167]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_168_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[168]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[168]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_169_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[169]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[169]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_170_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[170]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[170]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_171_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[171]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[171]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_172_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[172]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[172]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_173_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[173]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[173]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_174_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[174]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[174]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_175_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[175]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[175]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_176_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[176]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[176]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_177_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[177]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[177]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_178_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[178]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[178]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_179_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[179]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[179]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_180_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[180]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[180]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_181_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[181]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[181]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_182_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[182]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[182]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_183_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[183]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[183]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_184_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[184]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[184]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_185_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[185]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[185]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_186_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[186]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[186]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_187_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[187]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[187]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_188_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[188]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[188]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_189_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[189]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[189]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_190_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[190]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[190]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_191_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[191]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[191]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_192_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[192]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[192]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_193_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[193]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[193]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_194_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[194]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[194]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_195_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[195]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[195]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_196_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[196]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[196]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_197_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[197]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[197]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_198_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[198]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[198]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_199_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[199]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[199]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_200_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[200]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[200]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_201_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[201]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[201]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_202_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[202]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[202]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_203_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[203]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[203]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_204_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[204]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[204]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_205_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[205]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[205]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_206_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[206]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[206]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_207_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[207]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[207]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_208_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[208]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[208]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_209_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[209]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[209]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_210_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[210]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[210]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_211_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[211]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[211]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_212_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[212]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[212]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_213_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[213]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[213]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_214_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[214]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[214]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_215_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[215]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[215]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_216_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[216]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[216]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_217_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[217]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[217]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_218_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[218]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[218]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_219_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[219]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[219]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_220_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[220]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[220]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_221_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[221]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[221]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_222_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[222]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[222]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_223_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[223]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[223]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_224_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[224]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[224]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_225_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[225]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[225]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_226_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[226]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[226]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_227_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[227]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[227]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_228_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[228]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[228]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_229_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[229]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[229]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_230_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[230]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[230]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_231_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[231]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[231]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_232_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[232]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[232]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_233_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[233]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[233]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_234_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[234]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[234]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_235_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[235]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[235]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_236_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[236]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[236]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_237_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[237]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[237]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_238_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[238]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[238]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_239_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[239]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[239]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_240_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[240]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[240]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_241_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[241]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[241]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_242_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[242]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[242]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_243_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[243]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[243]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_244_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[244]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[244]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_245_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[245]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[245]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_246_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[246]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[246]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_247_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[247]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[247]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_248_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[248]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[248]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_249_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[249]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[249]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_250_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[250]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[250]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_251_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[251]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[251]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_252_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[252]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[252]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_253_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[253]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[253]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_254_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[254]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[254]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_din_q0_255_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_din_q0[255]), .I0(PE_wrapper297_U0_fifo_w_out_V_V_din_pass_0[255]) );
  assign PE_wrapper297_U0_fifo_w_out_V_V_din_pass_1 = PE_wrapper297_U0_fifo_w_out_V_V_din_q0;
  wire  fifo_w_PE_12_4_V_V_full_n_q0;
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) fifo_w_PE_12_4_V_V_full_n_q0_lut ( .O(fifo_w_PE_12_4_V_V_full_n_q0), .I0(fifo_w_PE_12_4_V_V_full_n_pass_1) );
  assign fifo_w_PE_12_4_V_V_full_n_pass_0 = fifo_w_PE_12_4_V_V_full_n_q0;
  wire  PE_wrapper297_U0_fifo_w_out_V_V_write_q0;
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper297_U0_fifo_w_out_V_V_write_q0_lut ( .O(PE_wrapper297_U0_fifo_w_out_V_V_write_q0), .I0(PE_wrapper297_U0_fifo_w_out_V_V_write_pass_0) );
  assign PE_wrapper297_U0_fifo_w_out_V_V_write_pass_1 = PE_wrapper297_U0_fifo_w_out_V_V_write_q0;
  wire [255:0] PE_wrapper310_U0_fifo_cin_out_V_V_din_q0;
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_0_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[0]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[0]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_1_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[1]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[1]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_2_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[2]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[2]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_3_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[3]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[3]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_4_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[4]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[4]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_5_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[5]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[5]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_6_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[6]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[6]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_7_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[7]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[7]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_8_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[8]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[8]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_9_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[9]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[9]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_10_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[10]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[10]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_11_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[11]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[11]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_12_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[12]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[12]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_13_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[13]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[13]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_14_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[14]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[14]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_15_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[15]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[15]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_16_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[16]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[16]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_17_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[17]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[17]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_18_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[18]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[18]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_19_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[19]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[19]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_20_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[20]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[20]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_21_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[21]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[21]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_22_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[22]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[22]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_23_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[23]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[23]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_24_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[24]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[24]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_25_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[25]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[25]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_26_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[26]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[26]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_27_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[27]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[27]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_28_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[28]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[28]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_29_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[29]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[29]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_30_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[30]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[30]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_31_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[31]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[31]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_32_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[32]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[32]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_33_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[33]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[33]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_34_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[34]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[34]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_35_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[35]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[35]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_36_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[36]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[36]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_37_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[37]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[37]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_38_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[38]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[38]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_39_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[39]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[39]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_40_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[40]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[40]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_41_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[41]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[41]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_42_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[42]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[42]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_43_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[43]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[43]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_44_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[44]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[44]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_45_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[45]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[45]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_46_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[46]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[46]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_47_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[47]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[47]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_48_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[48]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[48]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_49_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[49]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[49]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_50_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[50]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[50]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_51_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[51]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[51]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_52_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[52]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[52]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_53_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[53]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[53]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_54_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[54]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[54]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_55_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[55]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[55]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_56_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[56]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[56]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_57_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[57]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[57]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_58_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[58]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[58]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_59_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[59]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[59]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_60_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[60]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[60]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_61_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[61]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[61]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_62_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[62]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[62]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_63_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[63]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[63]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_64_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[64]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[64]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_65_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[65]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[65]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_66_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[66]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[66]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_67_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[67]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[67]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_68_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[68]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[68]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_69_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[69]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[69]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_70_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[70]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[70]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_71_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[71]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[71]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_72_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[72]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[72]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_73_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[73]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[73]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_74_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[74]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[74]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_75_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[75]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[75]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_76_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[76]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[76]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_77_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[77]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[77]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_78_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[78]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[78]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_79_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[79]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[79]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_80_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[80]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[80]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_81_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[81]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[81]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_82_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[82]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[82]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_83_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[83]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[83]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_84_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[84]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[84]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_85_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[85]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[85]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_86_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[86]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[86]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_87_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[87]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[87]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_88_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[88]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[88]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_89_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[89]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[89]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_90_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[90]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[90]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_91_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[91]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[91]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_92_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[92]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[92]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_93_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[93]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[93]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_94_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[94]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[94]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_95_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[95]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[95]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_96_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[96]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[96]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_97_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[97]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[97]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_98_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[98]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[98]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_99_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[99]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[99]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_100_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[100]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[100]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_101_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[101]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[101]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_102_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[102]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[102]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_103_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[103]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[103]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_104_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[104]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[104]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_105_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[105]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[105]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_106_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[106]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[106]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_107_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[107]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[107]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_108_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[108]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[108]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_109_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[109]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[109]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_110_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[110]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[110]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_111_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[111]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[111]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_112_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[112]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[112]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_113_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[113]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[113]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_114_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[114]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[114]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_115_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[115]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[115]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_116_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[116]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[116]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_117_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[117]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[117]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_118_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[118]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[118]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_119_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[119]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[119]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_120_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[120]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[120]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_121_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[121]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[121]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_122_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[122]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[122]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_123_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[123]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[123]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_124_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[124]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[124]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_125_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[125]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[125]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_126_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[126]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[126]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_127_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[127]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[127]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_128_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[128]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[128]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_129_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[129]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[129]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_130_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[130]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[130]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_131_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[131]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[131]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_132_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[132]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[132]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_133_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[133]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[133]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_134_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[134]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[134]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_135_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[135]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[135]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_136_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[136]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[136]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_137_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[137]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[137]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_138_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[138]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[138]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_139_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[139]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[139]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_140_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[140]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[140]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_141_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[141]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[141]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_142_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[142]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[142]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_143_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[143]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[143]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_144_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[144]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[144]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_145_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[145]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[145]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_146_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[146]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[146]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_147_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[147]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[147]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_148_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[148]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[148]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_149_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[149]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[149]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_150_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[150]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[150]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_151_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[151]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[151]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_152_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[152]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[152]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_153_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[153]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[153]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_154_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[154]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[154]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_155_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[155]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[155]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_156_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[156]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[156]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_157_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[157]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[157]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_158_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[158]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[158]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_159_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[159]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[159]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_160_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[160]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[160]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_161_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[161]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[161]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_162_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[162]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[162]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_163_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[163]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[163]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_164_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[164]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[164]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_165_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[165]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[165]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_166_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[166]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[166]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_167_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[167]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[167]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_168_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[168]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[168]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_169_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[169]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[169]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_170_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[170]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[170]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_171_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[171]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[171]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_172_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[172]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[172]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_173_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[173]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[173]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_174_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[174]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[174]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_175_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[175]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[175]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_176_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[176]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[176]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_177_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[177]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[177]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_178_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[178]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[178]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_179_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[179]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[179]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_180_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[180]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[180]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_181_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[181]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[181]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_182_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[182]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[182]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_183_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[183]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[183]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_184_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[184]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[184]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_185_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[185]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[185]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_186_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[186]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[186]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_187_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[187]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[187]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_188_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[188]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[188]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_189_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[189]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[189]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_190_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[190]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[190]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_191_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[191]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[191]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_192_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[192]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[192]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_193_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[193]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[193]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_194_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[194]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[194]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_195_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[195]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[195]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_196_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[196]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[196]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_197_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[197]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[197]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_198_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[198]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[198]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_199_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[199]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[199]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_200_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[200]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[200]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_201_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[201]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[201]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_202_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[202]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[202]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_203_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[203]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[203]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_204_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[204]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[204]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_205_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[205]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[205]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_206_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[206]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[206]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_207_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[207]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[207]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_208_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[208]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[208]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_209_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[209]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[209]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_210_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[210]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[210]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_211_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[211]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[211]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_212_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[212]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[212]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_213_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[213]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[213]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_214_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[214]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[214]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_215_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[215]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[215]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_216_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[216]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[216]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_217_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[217]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[217]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_218_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[218]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[218]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_219_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[219]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[219]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_220_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[220]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[220]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_221_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[221]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[221]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_222_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[222]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[222]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_223_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[223]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[223]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_224_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[224]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[224]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_225_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[225]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[225]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_226_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[226]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[226]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_227_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[227]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[227]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_228_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[228]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[228]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_229_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[229]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[229]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_230_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[230]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[230]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_231_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[231]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[231]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_232_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[232]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[232]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_233_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[233]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[233]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_234_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[234]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[234]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_235_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[235]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[235]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_236_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[236]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[236]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_237_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[237]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[237]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_238_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[238]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[238]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_239_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[239]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[239]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_240_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[240]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[240]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_241_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[241]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[241]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_242_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[242]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[242]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_243_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[243]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[243]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_244_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[244]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[244]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_245_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[245]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[245]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_246_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[246]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[246]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_247_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[247]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[247]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_248_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[248]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[248]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_249_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[249]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[249]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_250_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[250]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[250]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_251_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[251]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[251]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_252_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[252]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[252]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_253_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[253]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[253]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_254_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[254]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[254]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_din_q0_255_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_din_q0[255]), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_0[255]) );
  assign PE_wrapper310_U0_fifo_cin_out_V_V_din_pass_1 = PE_wrapper310_U0_fifo_cin_out_V_V_din_q0;
  wire  fifo_cin_PE_14_4_V_V_full_n_q0;
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) fifo_cin_PE_14_4_V_V_full_n_q0_lut ( .O(fifo_cin_PE_14_4_V_V_full_n_q0), .I0(fifo_cin_PE_14_4_V_V_full_n_pass_1) );
  assign fifo_cin_PE_14_4_V_V_full_n_pass_0 = fifo_cin_PE_14_4_V_V_full_n_q0;
  wire  PE_wrapper310_U0_fifo_cin_out_V_V_write_q0;
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper310_U0_fifo_cin_out_V_V_write_q0_lut ( .O(PE_wrapper310_U0_fifo_cin_out_V_V_write_q0), .I0(PE_wrapper310_U0_fifo_cin_out_V_V_write_pass_0) );
  assign PE_wrapper310_U0_fifo_cin_out_V_V_write_pass_1 = PE_wrapper310_U0_fifo_cin_out_V_V_write_q0;
  wire [255:0] PE_wrapper307_U0_fifo_cin_out_V_V_din_q0;
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_0_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[0]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[0]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_1_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[1]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[1]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_2_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[2]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[2]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_3_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[3]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[3]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_4_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[4]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[4]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_5_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[5]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[5]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_6_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[6]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[6]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_7_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[7]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[7]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_8_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[8]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[8]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_9_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[9]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[9]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_10_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[10]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[10]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_11_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[11]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[11]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_12_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[12]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[12]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_13_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[13]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[13]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_14_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[14]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[14]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_15_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[15]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[15]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_16_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[16]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[16]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_17_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[17]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[17]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_18_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[18]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[18]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_19_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[19]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[19]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_20_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[20]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[20]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_21_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[21]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[21]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_22_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[22]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[22]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_23_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[23]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[23]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_24_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[24]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[24]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_25_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[25]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[25]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_26_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[26]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[26]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_27_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[27]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[27]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_28_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[28]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[28]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_29_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[29]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[29]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_30_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[30]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[30]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_31_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[31]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[31]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_32_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[32]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[32]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_33_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[33]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[33]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_34_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[34]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[34]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_35_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[35]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[35]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_36_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[36]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[36]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_37_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[37]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[37]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_38_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[38]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[38]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_39_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[39]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[39]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_40_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[40]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[40]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_41_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[41]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[41]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_42_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[42]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[42]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_43_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[43]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[43]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_44_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[44]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[44]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_45_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[45]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[45]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_46_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[46]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[46]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_47_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[47]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[47]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_48_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[48]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[48]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_49_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[49]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[49]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_50_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[50]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[50]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_51_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[51]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[51]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_52_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[52]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[52]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_53_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[53]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[53]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_54_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[54]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[54]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_55_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[55]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[55]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_56_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[56]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[56]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_57_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[57]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[57]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_58_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[58]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[58]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_59_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[59]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[59]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_60_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[60]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[60]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_61_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[61]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[61]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_62_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[62]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[62]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_63_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[63]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[63]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_64_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[64]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[64]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_65_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[65]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[65]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_66_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[66]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[66]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_67_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[67]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[67]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_68_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[68]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[68]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_69_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[69]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[69]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_70_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[70]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[70]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_71_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[71]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[71]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_72_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[72]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[72]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_73_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[73]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[73]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_74_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[74]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[74]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_75_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[75]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[75]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_76_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[76]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[76]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_77_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[77]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[77]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_78_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[78]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[78]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_79_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[79]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[79]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_80_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[80]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[80]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_81_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[81]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[81]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_82_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[82]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[82]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_83_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[83]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[83]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_84_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[84]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[84]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_85_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[85]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[85]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_86_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[86]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[86]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_87_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[87]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[87]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_88_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[88]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[88]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_89_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[89]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[89]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_90_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[90]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[90]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_91_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[91]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[91]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_92_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[92]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[92]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_93_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[93]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[93]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_94_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[94]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[94]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_95_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[95]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[95]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_96_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[96]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[96]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_97_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[97]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[97]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_98_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[98]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[98]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_99_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[99]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[99]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_100_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[100]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[100]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_101_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[101]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[101]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_102_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[102]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[102]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_103_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[103]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[103]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_104_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[104]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[104]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_105_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[105]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[105]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_106_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[106]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[106]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_107_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[107]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[107]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_108_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[108]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[108]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_109_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[109]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[109]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_110_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[110]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[110]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_111_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[111]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[111]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_112_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[112]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[112]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_113_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[113]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[113]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_114_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[114]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[114]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_115_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[115]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[115]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_116_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[116]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[116]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_117_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[117]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[117]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_118_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[118]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[118]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_119_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[119]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[119]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_120_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[120]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[120]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_121_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[121]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[121]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_122_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[122]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[122]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_123_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[123]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[123]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_124_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[124]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[124]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_125_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[125]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[125]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_126_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[126]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[126]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_127_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[127]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[127]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_128_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[128]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[128]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_129_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[129]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[129]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_130_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[130]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[130]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_131_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[131]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[131]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_132_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[132]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[132]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_133_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[133]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[133]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_134_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[134]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[134]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_135_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[135]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[135]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_136_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[136]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[136]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_137_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[137]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[137]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_138_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[138]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[138]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_139_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[139]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[139]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_140_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[140]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[140]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_141_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[141]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[141]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_142_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[142]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[142]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_143_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[143]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[143]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_144_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[144]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[144]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_145_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[145]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[145]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_146_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[146]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[146]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_147_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[147]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[147]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_148_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[148]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[148]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_149_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[149]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[149]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_150_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[150]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[150]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_151_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[151]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[151]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_152_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[152]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[152]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_153_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[153]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[153]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_154_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[154]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[154]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_155_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[155]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[155]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_156_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[156]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[156]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_157_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[157]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[157]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_158_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[158]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[158]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_159_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[159]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[159]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_160_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[160]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[160]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_161_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[161]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[161]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_162_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[162]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[162]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_163_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[163]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[163]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_164_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[164]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[164]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_165_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[165]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[165]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_166_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[166]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[166]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_167_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[167]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[167]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_168_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[168]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[168]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_169_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[169]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[169]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_170_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[170]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[170]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_171_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[171]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[171]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_172_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[172]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[172]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_173_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[173]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[173]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_174_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[174]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[174]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_175_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[175]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[175]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_176_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[176]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[176]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_177_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[177]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[177]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_178_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[178]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[178]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_179_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[179]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[179]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_180_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[180]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[180]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_181_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[181]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[181]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_182_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[182]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[182]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_183_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[183]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[183]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_184_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[184]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[184]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_185_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[185]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[185]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_186_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[186]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[186]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_187_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[187]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[187]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_188_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[188]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[188]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_189_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[189]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[189]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_190_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[190]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[190]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_191_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[191]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[191]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_192_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[192]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[192]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_193_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[193]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[193]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_194_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[194]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[194]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_195_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[195]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[195]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_196_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[196]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[196]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_197_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[197]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[197]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_198_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[198]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[198]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_199_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[199]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[199]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_200_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[200]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[200]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_201_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[201]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[201]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_202_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[202]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[202]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_203_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[203]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[203]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_204_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[204]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[204]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_205_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[205]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[205]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_206_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[206]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[206]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_207_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[207]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[207]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_208_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[208]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[208]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_209_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[209]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[209]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_210_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[210]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[210]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_211_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[211]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[211]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_212_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[212]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[212]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_213_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[213]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[213]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_214_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[214]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[214]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_215_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[215]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[215]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_216_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[216]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[216]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_217_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[217]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[217]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_218_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[218]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[218]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_219_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[219]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[219]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_220_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[220]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[220]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_221_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[221]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[221]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_222_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[222]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[222]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_223_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[223]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[223]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_224_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[224]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[224]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_225_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[225]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[225]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_226_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[226]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[226]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_227_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[227]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[227]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_228_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[228]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[228]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_229_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[229]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[229]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_230_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[230]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[230]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_231_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[231]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[231]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_232_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[232]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[232]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_233_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[233]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[233]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_234_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[234]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[234]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_235_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[235]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[235]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_236_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[236]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[236]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_237_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[237]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[237]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_238_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[238]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[238]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_239_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[239]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[239]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_240_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[240]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[240]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_241_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[241]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[241]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_242_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[242]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[242]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_243_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[243]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[243]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_244_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[244]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[244]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_245_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[245]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[245]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_246_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[246]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[246]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_247_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[247]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[247]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_248_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[248]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[248]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_249_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[249]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[249]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_250_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[250]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[250]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_251_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[251]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[251]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_252_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[252]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[252]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_253_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[253]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[253]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_254_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[254]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[254]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_din_q0_255_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_din_q0[255]), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_0[255]) );
  assign PE_wrapper307_U0_fifo_cin_out_V_V_din_pass_1 = PE_wrapper307_U0_fifo_cin_out_V_V_din_q0;
  wire  fifo_cin_PE_14_1_V_V_full_n_q0;
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) fifo_cin_PE_14_1_V_V_full_n_q0_lut ( .O(fifo_cin_PE_14_1_V_V_full_n_q0), .I0(fifo_cin_PE_14_1_V_V_full_n_pass_1) );
  assign fifo_cin_PE_14_1_V_V_full_n_pass_0 = fifo_cin_PE_14_1_V_V_full_n_q0;
  wire  PE_wrapper307_U0_fifo_cin_out_V_V_write_q0;
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper307_U0_fifo_cin_out_V_V_write_q0_lut ( .O(PE_wrapper307_U0_fifo_cin_out_V_V_write_q0), .I0(PE_wrapper307_U0_fifo_cin_out_V_V_write_pass_0) );
  assign PE_wrapper307_U0_fifo_cin_out_V_V_write_pass_1 = PE_wrapper307_U0_fifo_cin_out_V_V_write_q0;
  wire [255:0] PE_wrapper250_U0_fifo_w_out_V_V_din_q0;
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_0_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[0]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[0]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_1_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[1]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[1]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_2_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[2]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[2]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_3_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[3]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[3]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_4_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[4]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[4]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_5_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[5]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[5]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_6_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[6]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[6]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_7_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[7]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[7]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_8_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[8]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[8]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_9_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[9]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[9]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_10_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[10]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[10]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_11_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[11]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[11]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_12_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[12]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[12]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_13_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[13]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[13]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_14_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[14]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[14]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_15_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[15]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[15]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_16_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[16]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[16]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_17_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[17]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[17]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_18_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[18]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[18]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_19_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[19]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[19]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_20_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[20]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[20]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_21_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[21]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[21]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_22_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[22]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[22]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_23_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[23]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[23]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_24_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[24]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[24]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_25_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[25]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[25]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_26_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[26]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[26]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_27_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[27]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[27]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_28_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[28]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[28]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_29_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[29]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[29]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_30_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[30]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[30]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_31_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[31]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[31]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_32_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[32]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[32]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_33_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[33]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[33]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_34_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[34]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[34]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_35_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[35]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[35]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_36_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[36]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[36]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_37_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[37]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[37]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_38_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[38]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[38]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_39_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[39]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[39]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_40_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[40]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[40]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_41_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[41]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[41]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_42_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[42]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[42]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_43_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[43]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[43]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_44_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[44]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[44]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_45_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[45]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[45]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_46_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[46]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[46]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_47_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[47]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[47]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_48_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[48]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[48]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_49_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[49]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[49]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_50_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[50]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[50]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_51_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[51]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[51]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_52_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[52]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[52]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_53_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[53]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[53]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_54_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[54]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[54]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_55_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[55]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[55]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_56_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[56]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[56]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_57_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[57]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[57]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_58_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[58]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[58]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_59_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[59]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[59]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_60_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[60]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[60]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_61_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[61]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[61]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_62_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[62]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[62]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_63_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[63]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[63]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_64_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[64]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[64]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_65_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[65]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[65]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_66_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[66]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[66]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_67_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[67]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[67]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_68_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[68]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[68]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_69_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[69]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[69]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_70_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[70]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[70]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_71_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[71]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[71]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_72_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[72]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[72]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_73_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[73]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[73]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_74_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[74]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[74]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_75_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[75]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[75]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_76_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[76]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[76]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_77_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[77]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[77]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_78_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[78]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[78]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_79_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[79]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[79]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_80_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[80]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[80]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_81_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[81]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[81]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_82_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[82]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[82]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_83_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[83]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[83]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_84_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[84]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[84]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_85_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[85]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[85]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_86_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[86]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[86]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_87_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[87]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[87]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_88_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[88]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[88]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_89_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[89]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[89]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_90_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[90]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[90]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_91_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[91]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[91]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_92_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[92]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[92]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_93_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[93]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[93]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_94_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[94]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[94]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_95_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[95]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[95]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_96_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[96]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[96]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_97_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[97]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[97]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_98_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[98]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[98]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_99_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[99]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[99]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_100_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[100]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[100]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_101_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[101]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[101]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_102_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[102]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[102]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_103_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[103]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[103]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_104_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[104]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[104]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_105_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[105]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[105]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_106_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[106]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[106]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_107_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[107]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[107]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_108_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[108]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[108]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_109_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[109]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[109]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_110_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[110]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[110]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_111_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[111]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[111]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_112_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[112]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[112]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_113_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[113]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[113]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_114_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[114]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[114]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_115_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[115]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[115]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_116_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[116]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[116]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_117_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[117]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[117]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_118_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[118]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[118]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_119_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[119]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[119]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_120_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[120]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[120]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_121_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[121]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[121]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_122_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[122]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[122]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_123_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[123]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[123]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_124_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[124]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[124]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_125_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[125]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[125]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_126_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[126]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[126]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_127_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[127]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[127]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_128_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[128]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[128]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_129_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[129]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[129]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_130_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[130]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[130]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_131_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[131]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[131]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_132_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[132]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[132]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_133_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[133]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[133]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_134_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[134]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[134]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_135_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[135]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[135]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_136_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[136]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[136]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_137_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[137]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[137]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_138_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[138]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[138]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_139_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[139]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[139]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_140_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[140]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[140]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_141_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[141]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[141]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_142_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[142]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[142]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_143_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[143]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[143]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_144_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[144]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[144]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_145_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[145]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[145]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_146_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[146]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[146]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_147_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[147]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[147]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_148_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[148]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[148]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_149_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[149]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[149]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_150_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[150]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[150]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_151_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[151]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[151]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_152_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[152]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[152]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_153_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[153]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[153]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_154_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[154]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[154]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_155_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[155]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[155]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_156_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[156]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[156]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_157_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[157]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[157]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_158_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[158]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[158]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_159_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[159]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[159]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_160_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[160]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[160]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_161_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[161]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[161]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_162_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[162]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[162]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_163_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[163]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[163]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_164_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[164]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[164]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_165_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[165]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[165]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_166_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[166]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[166]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_167_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[167]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[167]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_168_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[168]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[168]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_169_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[169]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[169]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_170_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[170]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[170]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_171_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[171]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[171]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_172_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[172]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[172]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_173_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[173]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[173]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_174_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[174]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[174]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_175_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[175]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[175]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_176_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[176]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[176]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_177_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[177]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[177]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_178_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[178]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[178]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_179_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[179]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[179]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_180_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[180]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[180]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_181_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[181]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[181]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_182_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[182]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[182]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_183_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[183]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[183]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_184_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[184]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[184]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_185_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[185]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[185]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_186_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[186]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[186]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_187_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[187]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[187]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_188_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[188]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[188]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_189_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[189]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[189]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_190_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[190]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[190]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_191_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[191]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[191]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_192_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[192]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[192]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_193_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[193]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[193]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_194_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[194]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[194]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_195_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[195]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[195]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_196_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[196]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[196]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_197_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[197]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[197]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_198_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[198]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[198]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_199_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[199]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[199]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_200_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[200]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[200]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_201_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[201]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[201]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_202_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[202]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[202]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_203_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[203]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[203]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_204_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[204]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[204]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_205_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[205]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[205]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_206_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[206]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[206]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_207_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[207]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[207]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_208_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[208]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[208]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_209_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[209]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[209]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_210_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[210]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[210]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_211_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[211]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[211]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_212_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[212]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[212]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_213_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[213]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[213]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_214_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[214]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[214]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_215_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[215]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[215]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_216_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[216]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[216]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_217_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[217]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[217]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_218_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[218]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[218]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_219_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[219]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[219]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_220_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[220]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[220]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_221_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[221]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[221]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_222_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[222]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[222]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_223_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[223]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[223]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_224_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[224]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[224]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_225_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[225]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[225]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_226_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[226]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[226]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_227_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[227]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[227]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_228_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[228]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[228]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_229_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[229]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[229]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_230_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[230]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[230]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_231_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[231]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[231]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_232_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[232]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[232]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_233_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[233]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[233]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_234_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[234]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[234]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_235_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[235]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[235]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_236_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[236]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[236]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_237_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[237]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[237]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_238_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[238]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[238]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_239_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[239]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[239]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_240_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[240]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[240]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_241_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[241]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[241]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_242_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[242]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[242]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_243_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[243]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[243]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_244_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[244]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[244]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_245_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[245]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[245]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_246_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[246]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[246]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_247_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[247]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[247]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_248_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[248]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[248]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_249_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[249]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[249]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_250_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[250]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[250]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_251_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[251]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[251]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_252_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[252]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[252]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_253_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[253]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[253]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_254_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[254]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[254]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_din_q0_255_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_din_q0[255]), .I0(PE_wrapper250_U0_fifo_w_out_V_V_din_pass_0[255]) );
  assign PE_wrapper250_U0_fifo_w_out_V_V_din_pass_1 = PE_wrapper250_U0_fifo_w_out_V_V_din_q0;
  wire  fifo_w_PE_8_5_V_V_full_n_q0;
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) fifo_w_PE_8_5_V_V_full_n_q0_lut ( .O(fifo_w_PE_8_5_V_V_full_n_q0), .I0(fifo_w_PE_8_5_V_V_full_n_pass_1) );
  assign fifo_w_PE_8_5_V_V_full_n_pass_0 = fifo_w_PE_8_5_V_V_full_n_q0;
  wire  PE_wrapper250_U0_fifo_w_out_V_V_write_q0;
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper250_U0_fifo_w_out_V_V_write_q0_lut ( .O(PE_wrapper250_U0_fifo_w_out_V_V_write_q0), .I0(PE_wrapper250_U0_fifo_w_out_V_V_write_pass_0) );
  assign PE_wrapper250_U0_fifo_w_out_V_V_write_pass_1 = PE_wrapper250_U0_fifo_w_out_V_V_write_q0;
  wire [255:0] PE_wrapper238_U0_fifo_w_out_V_V_din_q0;
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_0_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[0]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[0]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_1_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[1]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[1]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_2_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[2]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[2]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_3_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[3]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[3]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_4_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[4]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[4]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_5_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[5]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[5]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_6_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[6]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[6]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_7_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[7]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[7]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_8_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[8]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[8]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_9_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[9]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[9]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_10_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[10]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[10]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_11_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[11]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[11]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_12_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[12]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[12]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_13_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[13]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[13]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_14_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[14]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[14]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_15_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[15]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[15]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_16_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[16]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[16]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_17_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[17]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[17]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_18_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[18]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[18]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_19_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[19]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[19]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_20_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[20]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[20]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_21_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[21]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[21]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_22_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[22]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[22]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_23_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[23]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[23]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_24_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[24]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[24]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_25_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[25]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[25]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_26_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[26]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[26]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_27_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[27]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[27]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_28_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[28]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[28]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_29_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[29]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[29]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_30_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[30]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[30]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_31_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[31]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[31]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_32_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[32]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[32]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_33_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[33]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[33]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_34_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[34]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[34]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_35_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[35]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[35]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_36_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[36]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[36]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_37_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[37]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[37]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_38_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[38]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[38]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_39_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[39]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[39]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_40_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[40]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[40]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_41_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[41]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[41]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_42_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[42]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[42]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_43_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[43]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[43]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_44_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[44]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[44]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_45_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[45]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[45]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_46_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[46]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[46]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_47_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[47]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[47]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_48_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[48]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[48]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_49_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[49]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[49]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_50_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[50]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[50]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_51_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[51]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[51]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_52_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[52]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[52]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_53_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[53]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[53]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_54_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[54]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[54]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_55_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[55]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[55]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_56_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[56]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[56]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_57_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[57]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[57]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_58_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[58]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[58]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_59_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[59]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[59]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_60_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[60]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[60]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_61_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[61]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[61]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_62_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[62]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[62]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_63_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[63]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[63]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_64_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[64]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[64]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_65_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[65]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[65]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_66_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[66]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[66]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_67_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[67]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[67]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_68_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[68]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[68]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_69_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[69]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[69]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_70_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[70]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[70]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_71_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[71]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[71]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_72_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[72]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[72]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_73_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[73]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[73]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_74_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[74]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[74]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_75_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[75]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[75]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_76_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[76]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[76]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_77_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[77]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[77]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_78_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[78]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[78]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_79_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[79]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[79]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_80_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[80]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[80]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_81_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[81]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[81]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_82_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[82]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[82]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_83_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[83]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[83]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_84_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[84]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[84]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_85_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[85]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[85]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_86_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[86]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[86]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_87_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[87]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[87]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_88_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[88]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[88]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_89_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[89]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[89]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_90_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[90]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[90]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_91_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[91]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[91]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_92_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[92]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[92]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_93_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[93]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[93]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_94_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[94]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[94]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_95_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[95]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[95]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_96_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[96]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[96]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_97_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[97]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[97]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_98_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[98]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[98]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_99_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[99]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[99]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_100_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[100]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[100]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_101_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[101]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[101]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_102_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[102]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[102]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_103_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[103]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[103]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_104_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[104]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[104]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_105_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[105]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[105]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_106_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[106]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[106]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_107_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[107]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[107]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_108_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[108]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[108]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_109_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[109]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[109]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_110_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[110]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[110]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_111_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[111]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[111]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_112_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[112]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[112]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_113_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[113]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[113]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_114_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[114]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[114]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_115_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[115]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[115]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_116_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[116]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[116]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_117_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[117]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[117]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_118_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[118]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[118]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_119_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[119]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[119]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_120_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[120]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[120]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_121_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[121]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[121]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_122_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[122]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[122]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_123_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[123]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[123]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_124_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[124]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[124]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_125_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[125]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[125]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_126_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[126]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[126]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_127_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[127]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[127]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_128_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[128]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[128]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_129_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[129]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[129]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_130_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[130]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[130]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_131_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[131]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[131]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_132_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[132]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[132]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_133_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[133]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[133]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_134_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[134]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[134]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_135_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[135]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[135]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_136_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[136]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[136]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_137_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[137]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[137]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_138_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[138]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[138]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_139_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[139]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[139]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_140_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[140]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[140]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_141_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[141]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[141]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_142_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[142]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[142]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_143_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[143]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[143]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_144_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[144]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[144]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_145_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[145]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[145]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_146_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[146]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[146]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_147_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[147]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[147]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_148_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[148]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[148]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_149_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[149]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[149]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_150_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[150]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[150]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_151_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[151]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[151]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_152_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[152]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[152]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_153_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[153]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[153]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_154_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[154]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[154]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_155_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[155]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[155]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_156_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[156]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[156]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_157_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[157]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[157]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_158_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[158]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[158]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_159_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[159]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[159]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_160_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[160]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[160]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_161_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[161]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[161]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_162_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[162]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[162]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_163_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[163]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[163]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_164_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[164]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[164]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_165_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[165]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[165]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_166_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[166]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[166]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_167_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[167]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[167]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_168_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[168]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[168]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_169_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[169]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[169]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_170_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[170]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[170]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_171_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[171]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[171]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_172_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[172]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[172]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_173_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[173]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[173]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_174_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[174]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[174]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_175_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[175]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[175]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_176_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[176]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[176]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_177_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[177]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[177]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_178_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[178]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[178]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_179_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[179]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[179]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_180_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[180]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[180]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_181_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[181]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[181]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_182_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[182]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[182]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_183_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[183]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[183]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_184_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[184]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[184]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_185_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[185]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[185]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_186_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[186]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[186]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_187_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[187]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[187]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_188_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[188]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[188]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_189_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[189]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[189]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_190_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[190]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[190]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_191_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[191]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[191]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_192_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[192]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[192]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_193_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[193]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[193]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_194_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[194]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[194]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_195_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[195]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[195]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_196_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[196]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[196]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_197_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[197]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[197]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_198_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[198]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[198]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_199_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[199]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[199]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_200_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[200]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[200]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_201_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[201]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[201]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_202_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[202]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[202]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_203_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[203]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[203]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_204_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[204]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[204]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_205_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[205]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[205]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_206_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[206]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[206]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_207_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[207]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[207]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_208_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[208]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[208]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_209_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[209]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[209]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_210_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[210]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[210]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_211_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[211]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[211]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_212_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[212]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[212]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_213_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[213]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[213]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_214_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[214]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[214]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_215_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[215]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[215]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_216_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[216]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[216]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_217_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[217]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[217]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_218_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[218]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[218]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_219_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[219]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[219]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_220_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[220]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[220]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_221_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[221]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[221]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_222_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[222]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[222]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_223_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[223]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[223]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_224_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[224]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[224]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_225_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[225]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[225]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_226_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[226]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[226]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_227_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[227]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[227]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_228_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[228]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[228]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_229_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[229]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[229]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_230_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[230]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[230]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_231_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[231]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[231]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_232_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[232]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[232]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_233_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[233]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[233]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_234_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[234]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[234]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_235_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[235]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[235]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_236_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[236]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[236]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_237_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[237]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[237]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_238_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[238]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[238]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_239_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[239]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[239]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_240_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[240]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[240]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_241_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[241]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[241]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_242_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[242]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[242]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_243_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[243]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[243]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_244_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[244]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[244]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_245_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[245]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[245]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_246_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[246]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[246]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_247_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[247]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[247]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_248_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[248]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[248]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_249_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[249]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[249]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_250_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[250]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[250]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_251_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[251]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[251]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_252_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[252]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[252]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_253_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[253]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[253]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_254_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[254]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[254]) );
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_din_q0_255_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_din_q0[255]), .I0(PE_wrapper238_U0_fifo_w_out_V_V_din_pass_0[255]) );
  assign PE_wrapper238_U0_fifo_w_out_V_V_din_pass_1 = PE_wrapper238_U0_fifo_w_out_V_V_din_q0;
  wire  fifo_w_PE_7_5_V_V_full_n_q0;
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) fifo_w_PE_7_5_V_V_full_n_q0_lut ( .O(fifo_w_PE_7_5_V_V_full_n_q0), .I0(fifo_w_PE_7_5_V_V_full_n_pass_1) );
  assign fifo_w_PE_7_5_V_V_full_n_pass_0 = fifo_w_PE_7_5_V_V_full_n_q0;
  wire  PE_wrapper238_U0_fifo_w_out_V_V_write_q0;
(* dont_touch = "yes" *) LUT1 #(.INIT(2'b10)) PE_wrapper238_U0_fifo_w_out_V_V_write_q0_lut ( .O(PE_wrapper238_U0_fifo_w_out_V_V_write_q0), .I0(PE_wrapper238_U0_fifo_w_out_V_V_write_pass_0) );
  assign PE_wrapper238_U0_fifo_w_out_V_V_write_pass_1 = PE_wrapper238_U0_fifo_w_out_V_V_write_q0;
wire [31:0] PE_wrapper320_U0_fifo_cout_drain_out_V_din;
assign PE_wrapper320_U0_fifo_cout_drain_out_V_din_pass_0 = PE_wrapper320_U0_fifo_cout_drain_out_V_din;
wire  fifo_cout_drain_PE_14_2_V_full_n;
reg  fifo_cout_drain_PE_14_2_V_full_n_q_for_broadcast;
always @ (posedge ap_clk) fifo_cout_drain_PE_14_2_V_full_n_q_for_broadcast <= fifo_cout_drain_PE_14_2_V_full_n_pass_0;
assign fifo_cout_drain_PE_14_2_V_full_n = fifo_cout_drain_PE_14_2_V_full_n_q_for_broadcast;
wire  PE_wrapper320_U0_fifo_cout_drain_out_V_write;
assign PE_wrapper320_U0_fifo_cout_drain_out_V_write_pass_0 = PE_wrapper320_U0_fifo_cout_drain_out_V_write;
wire [63:0] cout_drain_IO_L1_out_wrapper433_U0_fifo_cout_drain_out_V_V_din;
assign cout_drain_IO_L1_out_wrapper433_U0_fifo_cout_drain_out_V_V_din = cout_drain_IO_L1_out_wrapper433_U0_fifo_cout_drain_out_V_V_din_pass_0;
wire  fifo_cout_drain_cout_drain_IO_L1_out_4_13_V_V_full_n;
assign fifo_cout_drain_cout_drain_IO_L1_out_4_13_V_V_full_n_pass_0 = fifo_cout_drain_cout_drain_IO_L1_out_4_13_V_V_full_n;
wire  cout_drain_IO_L1_out_wrapper433_U0_fifo_cout_drain_out_V_V_write;
assign cout_drain_IO_L1_out_wrapper433_U0_fifo_cout_drain_out_V_V_write = cout_drain_IO_L1_out_wrapper433_U0_fifo_cout_drain_out_V_V_write_pass_0;
wire [255:0] PE_wrapper309_U0_fifo_cin_out_V_V_din;
assign PE_wrapper309_U0_fifo_cin_out_V_V_din = PE_wrapper309_U0_fifo_cin_out_V_V_din_pass_1;
wire  fifo_cin_PE_14_3_V_V_full_n;
assign fifo_cin_PE_14_3_V_V_full_n_pass_1 = fifo_cin_PE_14_3_V_V_full_n;
wire  PE_wrapper309_U0_fifo_cin_out_V_V_write;
assign PE_wrapper309_U0_fifo_cin_out_V_V_write = PE_wrapper309_U0_fifo_cin_out_V_V_write_pass_1;
wire [63:0] cout_drain_IO_L1_out_wrapper402_U0_fifo_cout_drain_out_V_V_din;
assign cout_drain_IO_L1_out_wrapper402_U0_fifo_cout_drain_out_V_V_din_pass_0 = cout_drain_IO_L1_out_wrapper402_U0_fifo_cout_drain_out_V_V_din;
wire  fifo_cout_drain_cout_drain_IO_L1_out_2_12_V_V_full_n;
reg  fifo_cout_drain_cout_drain_IO_L1_out_2_12_V_V_full_n_q_for_broadcast;
always @ (posedge ap_clk) fifo_cout_drain_cout_drain_IO_L1_out_2_12_V_V_full_n_q_for_broadcast <= fifo_cout_drain_cout_drain_IO_L1_out_2_12_V_V_full_n_pass_0;
assign fifo_cout_drain_cout_drain_IO_L1_out_2_12_V_V_full_n = fifo_cout_drain_cout_drain_IO_L1_out_2_12_V_V_full_n_q_for_broadcast;
wire  cout_drain_IO_L1_out_wrapper402_U0_fifo_cout_drain_out_V_V_write;
assign cout_drain_IO_L1_out_wrapper402_U0_fifo_cout_drain_out_V_V_write_pass_0 = cout_drain_IO_L1_out_wrapper402_U0_fifo_cout_drain_out_V_V_write;
wire [255:0] w_IO_L2_in149_U0_fifo_w_out_V_V_din;
assign w_IO_L2_in149_U0_fifo_w_out_V_V_din_pass_0 = w_IO_L2_in149_U0_fifo_w_out_V_V_din;
wire  fifo_w_w_IO_L2_in_15_V_V_full_n;
reg  fifo_w_w_IO_L2_in_15_V_V_full_n_q_for_broadcast;
always @ (posedge ap_clk) fifo_w_w_IO_L2_in_15_V_V_full_n_q_for_broadcast <= fifo_w_w_IO_L2_in_15_V_V_full_n_pass_0;
assign fifo_w_w_IO_L2_in_15_V_V_full_n = fifo_w_w_IO_L2_in_15_V_V_full_n_q_for_broadcast;
wire  w_IO_L2_in149_U0_fifo_w_out_V_V_write;
assign w_IO_L2_in149_U0_fifo_w_out_V_V_write_pass_0 = w_IO_L2_in149_U0_fifo_w_out_V_V_write;
wire [31:0] PE_wrapper286_U0_fifo_cout_drain_out_V_din;
assign PE_wrapper286_U0_fifo_cout_drain_out_V_din_pass_0 = PE_wrapper286_U0_fifo_cout_drain_out_V_din;
wire  fifo_cout_drain_PE_11_4_V_full_n;
reg  fifo_cout_drain_PE_11_4_V_full_n_q_for_broadcast;
always @ (posedge ap_clk) fifo_cout_drain_PE_11_4_V_full_n_q_for_broadcast <= fifo_cout_drain_PE_11_4_V_full_n_pass_0;
assign fifo_cout_drain_PE_11_4_V_full_n = fifo_cout_drain_PE_11_4_V_full_n_q_for_broadcast;
wire  PE_wrapper286_U0_fifo_cout_drain_out_V_write;
assign PE_wrapper286_U0_fifo_cout_drain_out_V_write_pass_0 = PE_wrapper286_U0_fifo_cout_drain_out_V_write;
wire [255:0] PE_wrapper214_U0_fifo_cin_out_V_V_din;
assign PE_wrapper214_U0_fifo_cin_out_V_V_din = PE_wrapper214_U0_fifo_cin_out_V_V_din_pass_1;
wire  fifo_cin_PE_6_4_V_V_full_n;
assign fifo_cin_PE_6_4_V_V_full_n_pass_1 = fifo_cin_PE_6_4_V_V_full_n;
wire  PE_wrapper214_U0_fifo_cin_out_V_V_write;
assign PE_wrapper214_U0_fifo_cin_out_V_V_write = PE_wrapper214_U0_fifo_cin_out_V_V_write_pass_1;
wire [63:0] cout_drain_IO_L1_out_wrapper432_U0_fifo_cout_drain_out_V_V_din;
assign cout_drain_IO_L1_out_wrapper432_U0_fifo_cout_drain_out_V_V_din_pass_0 = cout_drain_IO_L1_out_wrapper432_U0_fifo_cout_drain_out_V_V_din;
wire  fifo_cout_drain_cout_drain_IO_L1_out_4_14_V_V_full_n;
reg  fifo_cout_drain_cout_drain_IO_L1_out_4_14_V_V_full_n_q_for_broadcast;
always @ (posedge ap_clk) fifo_cout_drain_cout_drain_IO_L1_out_4_14_V_V_full_n_q_for_broadcast <= fifo_cout_drain_cout_drain_IO_L1_out_4_14_V_V_full_n_pass_0;
assign fifo_cout_drain_cout_drain_IO_L1_out_4_14_V_V_full_n = fifo_cout_drain_cout_drain_IO_L1_out_4_14_V_V_full_n_q_for_broadcast;
wire  cout_drain_IO_L1_out_wrapper432_U0_fifo_cout_drain_out_V_V_write;
assign cout_drain_IO_L1_out_wrapper432_U0_fifo_cout_drain_out_V_V_write_pass_0 = cout_drain_IO_L1_out_wrapper432_U0_fifo_cout_drain_out_V_V_write;
wire [255:0] PE_wrapper318_U0_fifo_w_out_V_V_din;
assign PE_wrapper318_U0_fifo_w_out_V_V_din_pass_0 = PE_wrapper318_U0_fifo_w_out_V_V_din;
wire  fifo_w_PE_14_1_V_V_full_n;
reg  fifo_w_PE_14_1_V_V_full_n_q_for_broadcast;
always @ (posedge ap_clk) fifo_w_PE_14_1_V_V_full_n_q_for_broadcast <= fifo_w_PE_14_1_V_V_full_n_pass_0;
assign fifo_w_PE_14_1_V_V_full_n = fifo_w_PE_14_1_V_V_full_n_q_for_broadcast;
wire  PE_wrapper318_U0_fifo_w_out_V_V_write;
assign PE_wrapper318_U0_fifo_w_out_V_V_write_pass_0 = PE_wrapper318_U0_fifo_w_out_V_V_write;
wire [31:0] PE_wrapper226_U0_fifo_cout_drain_out_V_din;
assign PE_wrapper226_U0_fifo_cout_drain_out_V_din_pass_0 = PE_wrapper226_U0_fifo_cout_drain_out_V_din;
wire  fifo_cout_drain_PE_6_4_V_full_n;
reg  fifo_cout_drain_PE_6_4_V_full_n_q_for_broadcast;
always @ (posedge ap_clk) fifo_cout_drain_PE_6_4_V_full_n_q_for_broadcast <= fifo_cout_drain_PE_6_4_V_full_n_pass_0;
assign fifo_cout_drain_PE_6_4_V_full_n = fifo_cout_drain_PE_6_4_V_full_n_q_for_broadcast;
wire  PE_wrapper226_U0_fifo_cout_drain_out_V_write;
assign PE_wrapper226_U0_fifo_cout_drain_out_V_write_pass_0 = PE_wrapper226_U0_fifo_cout_drain_out_V_write;
wire [255:0] PE_wrapper286_U0_fifo_cin_out_V_V_din;
assign PE_wrapper286_U0_fifo_cin_out_V_V_din_pass_0 = PE_wrapper286_U0_fifo_cin_out_V_V_din;
wire  fifo_cin_PE_12_4_V_V_full_n;
reg  fifo_cin_PE_12_4_V_V_full_n_q_for_broadcast;
always @ (posedge ap_clk) fifo_cin_PE_12_4_V_V_full_n_q_for_broadcast <= fifo_cin_PE_12_4_V_V_full_n_pass_0;
assign fifo_cin_PE_12_4_V_V_full_n = fifo_cin_PE_12_4_V_V_full_n_q_for_broadcast;
wire  PE_wrapper286_U0_fifo_cin_out_V_V_write;
assign PE_wrapper286_U0_fifo_cin_out_V_V_write_pass_0 = PE_wrapper286_U0_fifo_cin_out_V_V_write;
wire [255:0] w_IO_L2_in148_U0_fifo_w_out_V_V_din;
assign w_IO_L2_in148_U0_fifo_w_out_V_V_din = w_IO_L2_in148_U0_fifo_w_out_V_V_din_pass_0;
wire  fifo_w_w_IO_L2_in_14_V_V_full_n;
assign fifo_w_w_IO_L2_in_14_V_V_full_n_pass_0 = fifo_w_w_IO_L2_in_14_V_V_full_n;
wire  w_IO_L2_in148_U0_fifo_w_out_V_V_write;
assign w_IO_L2_in148_U0_fifo_w_out_V_V_write = w_IO_L2_in148_U0_fifo_w_out_V_V_write_pass_0;
wire [255:0] PE_wrapper320_U0_fifo_cin_out_V_V_din;
assign PE_wrapper320_U0_fifo_cin_out_V_V_din_pass_0 = PE_wrapper320_U0_fifo_cin_out_V_V_din;
wire  fifo_cin_PE_15_2_V_V_full_n;
reg  fifo_cin_PE_15_2_V_V_full_n_q_for_broadcast;
always @ (posedge ap_clk) fifo_cin_PE_15_2_V_V_full_n_q_for_broadcast <= fifo_cin_PE_15_2_V_V_full_n_pass_0;
assign fifo_cin_PE_15_2_V_V_full_n = fifo_cin_PE_15_2_V_V_full_n_q_for_broadcast;
wire  PE_wrapper320_U0_fifo_cin_out_V_V_write;
assign PE_wrapper320_U0_fifo_cin_out_V_V_write_pass_0 = PE_wrapper320_U0_fifo_cin_out_V_V_write;
wire [63:0] cout_drain_IO_L1_out_wrapper418_U0_fifo_cout_drain_out_V_V_din;
assign cout_drain_IO_L1_out_wrapper418_U0_fifo_cout_drain_out_V_V_din = cout_drain_IO_L1_out_wrapper418_U0_fifo_cout_drain_out_V_V_din_pass_1;
wire  fifo_cout_drain_cout_drain_IO_L1_out_3_12_V_V_full_n;
assign fifo_cout_drain_cout_drain_IO_L1_out_3_12_V_V_full_n_pass_1 = fifo_cout_drain_cout_drain_IO_L1_out_3_12_V_V_full_n;
wire  cout_drain_IO_L1_out_wrapper418_U0_fifo_cout_drain_out_V_V_write;
assign cout_drain_IO_L1_out_wrapper418_U0_fifo_cout_drain_out_V_V_write = cout_drain_IO_L1_out_wrapper418_U0_fifo_cout_drain_out_V_V_write_pass_1;
wire [255:0] PE_wrapper225_U0_fifo_w_out_V_V_din;
assign PE_wrapper225_U0_fifo_w_out_V_V_din = PE_wrapper225_U0_fifo_w_out_V_V_din_pass_1;
wire  fifo_w_PE_6_4_V_V_full_n;
assign fifo_w_PE_6_4_V_V_full_n_pass_1 = fifo_w_PE_6_4_V_V_full_n;
wire  PE_wrapper225_U0_fifo_w_out_V_V_write;
assign PE_wrapper225_U0_fifo_w_out_V_V_write = PE_wrapper225_U0_fifo_w_out_V_V_write_pass_1;
wire [63:0] cout_drain_IO_L1_out_wrapper416_U0_fifo_cout_drain_out_V_V_din;
assign cout_drain_IO_L1_out_wrapper416_U0_fifo_cout_drain_out_V_V_din_pass_0 = cout_drain_IO_L1_out_wrapper416_U0_fifo_cout_drain_out_V_V_din;
wire  fifo_cout_drain_cout_drain_IO_L1_out_3_14_V_V_full_n;
reg  fifo_cout_drain_cout_drain_IO_L1_out_3_14_V_V_full_n_q_for_broadcast;
always @ (posedge ap_clk) fifo_cout_drain_cout_drain_IO_L1_out_3_14_V_V_full_n_q_for_broadcast <= fifo_cout_drain_cout_drain_IO_L1_out_3_14_V_V_full_n_pass_0;
assign fifo_cout_drain_cout_drain_IO_L1_out_3_14_V_V_full_n = fifo_cout_drain_cout_drain_IO_L1_out_3_14_V_V_full_n_q_for_broadcast;
wire  cout_drain_IO_L1_out_wrapper416_U0_fifo_cout_drain_out_V_V_write;
assign cout_drain_IO_L1_out_wrapper416_U0_fifo_cout_drain_out_V_V_write_pass_0 = cout_drain_IO_L1_out_wrapper416_U0_fifo_cout_drain_out_V_V_write;
wire [255:0] PE_wrapper330_U0_fifo_cin_out_V_V_din;
assign PE_wrapper330_U0_fifo_cin_out_V_V_din_pass_0 = PE_wrapper330_U0_fifo_cin_out_V_V_din;
wire  fifo_cin_PE_16_0_V_V_full_n;
reg  fifo_cin_PE_16_0_V_V_full_n_q_for_broadcast;
always @ (posedge ap_clk) fifo_cin_PE_16_0_V_V_full_n_q_for_broadcast <= fifo_cin_PE_16_0_V_V_full_n_pass_0;
assign fifo_cin_PE_16_0_V_V_full_n = fifo_cin_PE_16_0_V_V_full_n_q_for_broadcast;
wire  PE_wrapper330_U0_fifo_cin_out_V_V_write;
assign PE_wrapper330_U0_fifo_cin_out_V_V_write_pass_0 = PE_wrapper330_U0_fifo_cin_out_V_V_write;
wire [255:0] PE_wrapper330_U0_fifo_w_out_V_V_din;
assign PE_wrapper330_U0_fifo_w_out_V_V_din_pass_0 = PE_wrapper330_U0_fifo_w_out_V_V_din;
wire  fifo_w_PE_15_1_V_V_full_n;
reg  fifo_w_PE_15_1_V_V_full_n_q_for_broadcast;
always @ (posedge ap_clk) fifo_w_PE_15_1_V_V_full_n_q_for_broadcast <= fifo_w_PE_15_1_V_V_full_n_pass_0;
assign fifo_w_PE_15_1_V_V_full_n = fifo_w_PE_15_1_V_V_full_n_q_for_broadcast;
wire  PE_wrapper330_U0_fifo_w_out_V_V_write;
assign PE_wrapper330_U0_fifo_w_out_V_V_write_pass_0 = PE_wrapper330_U0_fifo_w_out_V_V_write;
wire [255:0] PE_wrapper285_U0_fifo_w_out_V_V_din;
assign PE_wrapper285_U0_fifo_w_out_V_V_din = PE_wrapper285_U0_fifo_w_out_V_V_din_pass_1;
wire  fifo_w_PE_11_4_V_V_full_n;
assign fifo_w_PE_11_4_V_V_full_n_pass_1 = fifo_w_PE_11_4_V_V_full_n;
wire  PE_wrapper285_U0_fifo_w_out_V_V_write;
assign PE_wrapper285_U0_fifo_w_out_V_V_write = PE_wrapper285_U0_fifo_w_out_V_V_write_pass_1;
wire [63:0] cout_drain_IO_L1_out_wrapper419_U0_fifo_cout_drain_out_V_V_din;
assign cout_drain_IO_L1_out_wrapper419_U0_fifo_cout_drain_out_V_V_din_pass_0 = cout_drain_IO_L1_out_wrapper419_U0_fifo_cout_drain_out_V_V_din;
wire  fifo_cout_drain_cout_drain_IO_L1_out_3_11_V_V_full_n;
reg  fifo_cout_drain_cout_drain_IO_L1_out_3_11_V_V_full_n_q_for_broadcast;
always @ (posedge ap_clk) fifo_cout_drain_cout_drain_IO_L1_out_3_11_V_V_full_n_q_for_broadcast <= fifo_cout_drain_cout_drain_IO_L1_out_3_11_V_V_full_n_pass_0;
assign fifo_cout_drain_cout_drain_IO_L1_out_3_11_V_V_full_n = fifo_cout_drain_cout_drain_IO_L1_out_3_11_V_V_full_n_q_for_broadcast;
wire  cout_drain_IO_L1_out_wrapper419_U0_fifo_cout_drain_out_V_V_write;
assign cout_drain_IO_L1_out_wrapper419_U0_fifo_cout_drain_out_V_V_write_pass_0 = cout_drain_IO_L1_out_wrapper419_U0_fifo_cout_drain_out_V_V_write;
wire [255:0] w_IO_L2_in_boundary_U0_fifo_w_local_out_V_V_din;
assign w_IO_L2_in_boundary_U0_fifo_w_local_out_V_V_din = w_IO_L2_in_boundary_U0_fifo_w_local_out_V_V_din_pass_0;
wire  fifo_w_PE_15_0_V_V_full_n;
assign fifo_w_PE_15_0_V_V_full_n_pass_0 = fifo_w_PE_15_0_V_V_full_n;
wire  w_IO_L2_in_boundary_U0_fifo_w_local_out_V_V_write;
assign w_IO_L2_in_boundary_U0_fifo_w_local_out_V_V_write = w_IO_L2_in_boundary_U0_fifo_w_local_out_V_V_write_pass_0;
wire [255:0] PE_wrapper273_U0_fifo_w_out_V_V_din;
assign PE_wrapper273_U0_fifo_w_out_V_V_din = PE_wrapper273_U0_fifo_w_out_V_V_din_pass_0;
wire  fifo_w_PE_10_4_V_V_full_n;
assign fifo_w_PE_10_4_V_V_full_n_pass_0 = fifo_w_PE_10_4_V_V_full_n;
wire  PE_wrapper273_U0_fifo_w_out_V_V_write;
assign PE_wrapper273_U0_fifo_w_out_V_V_write = PE_wrapper273_U0_fifo_w_out_V_V_write_pass_0;
wire [255:0] PE_wrapper286_U0_fifo_w_out_V_V_din;
assign PE_wrapper286_U0_fifo_w_out_V_V_din_pass_0 = PE_wrapper286_U0_fifo_w_out_V_V_din;
wire  fifo_w_PE_11_5_V_V_full_n;
reg  fifo_w_PE_11_5_V_V_full_n_q_for_broadcast;
always @ (posedge ap_clk) fifo_w_PE_11_5_V_V_full_n_q_for_broadcast <= fifo_w_PE_11_5_V_V_full_n_pass_0;
assign fifo_w_PE_11_5_V_V_full_n = fifo_w_PE_11_5_V_V_full_n_q_for_broadcast;
wire  PE_wrapper286_U0_fifo_w_out_V_V_write;
assign PE_wrapper286_U0_fifo_w_out_V_V_write_pass_0 = PE_wrapper286_U0_fifo_w_out_V_V_write;
wire [63:0] cout_drain_IO_L1_out_boundary_wrapper383_U0_fifo_cout_drain_out_V_V_din;
assign cout_drain_IO_L1_out_boundary_wrapper383_U0_fifo_cout_drain_out_V_V_din = cout_drain_IO_L1_out_boundary_wrapper383_U0_fifo_cout_drain_out_V_V_din_pass_0;
wire  fifo_cout_drain_cout_drain_IO_L1_out_1_15_V_V_full_n;
assign fifo_cout_drain_cout_drain_IO_L1_out_1_15_V_V_full_n_pass_0 = fifo_cout_drain_cout_drain_IO_L1_out_1_15_V_V_full_n;
wire  cout_drain_IO_L1_out_boundary_wrapper383_U0_fifo_cout_drain_out_V_V_write;
assign cout_drain_IO_L1_out_boundary_wrapper383_U0_fifo_cout_drain_out_V_V_write = cout_drain_IO_L1_out_boundary_wrapper383_U0_fifo_cout_drain_out_V_V_write_pass_0;
wire [31:0] PE_wrapper330_U0_fifo_cout_drain_out_V_din;
assign PE_wrapper330_U0_fifo_cout_drain_out_V_din_pass_0 = PE_wrapper330_U0_fifo_cout_drain_out_V_din;
wire  fifo_cout_drain_PE_15_0_V_full_n;
reg  fifo_cout_drain_PE_15_0_V_full_n_q_for_broadcast;
always @ (posedge ap_clk) fifo_cout_drain_PE_15_0_V_full_n_q_for_broadcast <= fifo_cout_drain_PE_15_0_V_full_n_pass_0;
assign fifo_cout_drain_PE_15_0_V_full_n = fifo_cout_drain_PE_15_0_V_full_n_q_for_broadcast;
wire  PE_wrapper330_U0_fifo_cout_drain_out_V_write;
assign PE_wrapper330_U0_fifo_cout_drain_out_V_write_pass_0 = PE_wrapper330_U0_fifo_cout_drain_out_V_write;
wire [255:0] PE_wrapper306_U0_fifo_cin_out_V_V_din;
assign PE_wrapper306_U0_fifo_cin_out_V_V_din = PE_wrapper306_U0_fifo_cin_out_V_V_din_pass_1;
wire  fifo_cin_PE_14_0_V_V_full_n;
assign fifo_cin_PE_14_0_V_V_full_n_pass_1 = fifo_cin_PE_14_0_V_V_full_n;
wire  PE_wrapper306_U0_fifo_cin_out_V_V_write;
assign PE_wrapper306_U0_fifo_cin_out_V_V_write = PE_wrapper306_U0_fifo_cin_out_V_V_write_pass_1;
wire [255:0] PE_wrapper321_U0_fifo_cin_out_V_V_din;
assign PE_wrapper321_U0_fifo_cin_out_V_V_din_pass_0 = PE_wrapper321_U0_fifo_cin_out_V_V_din;
wire  fifo_cin_PE_15_3_V_V_full_n;
reg  fifo_cin_PE_15_3_V_V_full_n_q_for_broadcast;
always @ (posedge ap_clk) fifo_cin_PE_15_3_V_V_full_n_q_for_broadcast <= fifo_cin_PE_15_3_V_V_full_n_pass_0;
assign fifo_cin_PE_15_3_V_V_full_n = fifo_cin_PE_15_3_V_V_full_n_q_for_broadcast;
wire  PE_wrapper321_U0_fifo_cin_out_V_V_write;
assign PE_wrapper321_U0_fifo_cin_out_V_V_write_pass_0 = PE_wrapper321_U0_fifo_cin_out_V_V_write;
wire [31:0] PE_wrapper285_U0_fifo_cout_drain_out_V_din;
assign PE_wrapper285_U0_fifo_cout_drain_out_V_din = PE_wrapper285_U0_fifo_cout_drain_out_V_din_pass_1;
wire  fifo_cout_drain_PE_11_3_V_full_n;
assign fifo_cout_drain_PE_11_3_V_full_n_pass_1 = fifo_cout_drain_PE_11_3_V_full_n;
wire  PE_wrapper285_U0_fifo_cout_drain_out_V_write;
assign PE_wrapper285_U0_fifo_cout_drain_out_V_write = PE_wrapper285_U0_fifo_cout_drain_out_V_write_pass_1;
wire [255:0] PE_wrapper319_U0_fifo_w_out_V_V_din;
assign PE_wrapper319_U0_fifo_w_out_V_V_din = PE_wrapper319_U0_fifo_w_out_V_V_din_pass_0;
wire  fifo_w_PE_14_2_V_V_full_n;
assign fifo_w_PE_14_2_V_V_full_n_pass_0 = fifo_w_PE_14_2_V_V_full_n;
wire  PE_wrapper319_U0_fifo_w_out_V_V_write;
assign PE_wrapper319_U0_fifo_w_out_V_V_write = PE_wrapper319_U0_fifo_w_out_V_V_write_pass_0;
wire [255:0] PE_wrapper226_U0_fifo_w_out_V_V_din;
assign PE_wrapper226_U0_fifo_w_out_V_V_din_pass_0 = PE_wrapper226_U0_fifo_w_out_V_V_din;
wire  fifo_w_PE_6_5_V_V_full_n;
reg  fifo_w_PE_6_5_V_V_full_n_q_for_broadcast;
always @ (posedge ap_clk) fifo_w_PE_6_5_V_V_full_n_q_for_broadcast <= fifo_w_PE_6_5_V_V_full_n_pass_0;
assign fifo_w_PE_6_5_V_V_full_n = fifo_w_PE_6_5_V_V_full_n_q_for_broadcast;
wire  PE_wrapper226_U0_fifo_w_out_V_V_write;
assign PE_wrapper226_U0_fifo_w_out_V_V_write_pass_0 = PE_wrapper226_U0_fifo_w_out_V_V_write;
wire [255:0] PE_wrapper308_U0_fifo_cin_out_V_V_din;
assign PE_wrapper308_U0_fifo_cin_out_V_V_din = PE_wrapper308_U0_fifo_cin_out_V_V_din_pass_0;
wire  fifo_cin_PE_14_2_V_V_full_n;
assign fifo_cin_PE_14_2_V_V_full_n_pass_0 = fifo_cin_PE_14_2_V_V_full_n;
wire  PE_wrapper308_U0_fifo_cin_out_V_V_write;
assign PE_wrapper308_U0_fifo_cin_out_V_V_write = PE_wrapper308_U0_fifo_cin_out_V_V_write_pass_0;
wire [63:0] cout_drain_IO_L1_out_wrapper384_U0_fifo_cout_drain_out_V_V_din;
assign cout_drain_IO_L1_out_wrapper384_U0_fifo_cout_drain_out_V_V_din_pass_0 = cout_drain_IO_L1_out_wrapper384_U0_fifo_cout_drain_out_V_V_din;
wire  fifo_cout_drain_cout_drain_IO_L1_out_1_14_V_V_full_n;
reg  fifo_cout_drain_cout_drain_IO_L1_out_1_14_V_V_full_n_q_for_broadcast;
always @ (posedge ap_clk) fifo_cout_drain_cout_drain_IO_L1_out_1_14_V_V_full_n_q_for_broadcast <= fifo_cout_drain_cout_drain_IO_L1_out_1_14_V_V_full_n_pass_0;
assign fifo_cout_drain_cout_drain_IO_L1_out_1_14_V_V_full_n = fifo_cout_drain_cout_drain_IO_L1_out_1_14_V_V_full_n_q_for_broadcast;
wire  cout_drain_IO_L1_out_wrapper384_U0_fifo_cout_drain_out_V_V_write;
assign cout_drain_IO_L1_out_wrapper384_U0_fifo_cout_drain_out_V_V_write_pass_0 = cout_drain_IO_L1_out_wrapper384_U0_fifo_cout_drain_out_V_V_write;
wire [31:0] PE_wrapper319_U0_fifo_cout_drain_out_V_din;
assign PE_wrapper319_U0_fifo_cout_drain_out_V_din = PE_wrapper319_U0_fifo_cout_drain_out_V_din_pass_0;
wire  fifo_cout_drain_PE_14_1_V_full_n;
assign fifo_cout_drain_PE_14_1_V_full_n_pass_0 = fifo_cout_drain_PE_14_1_V_full_n;
wire  PE_wrapper319_U0_fifo_cout_drain_out_V_write;
assign PE_wrapper319_U0_fifo_cout_drain_out_V_write = PE_wrapper319_U0_fifo_cout_drain_out_V_write_pass_0;
wire [31:0] PE_wrapper334_U0_fifo_cout_drain_out_V_din;
assign PE_wrapper334_U0_fifo_cout_drain_out_V_din = PE_wrapper334_U0_fifo_cout_drain_out_V_din_pass_0;
wire  fifo_cout_drain_PE_15_4_V_full_n;
assign fifo_cout_drain_PE_15_4_V_full_n_pass_0 = fifo_cout_drain_PE_15_4_V_full_n;
wire  PE_wrapper334_U0_fifo_cout_drain_out_V_write;
assign PE_wrapper334_U0_fifo_cout_drain_out_V_write = PE_wrapper334_U0_fifo_cout_drain_out_V_write_pass_0;
wire [63:0] cout_drain_IO_L1_out_boundary_wrapper415_U0_fifo_cout_drain_out_V_V_din;
assign cout_drain_IO_L1_out_boundary_wrapper415_U0_fifo_cout_drain_out_V_V_din = cout_drain_IO_L1_out_boundary_wrapper415_U0_fifo_cout_drain_out_V_V_din_pass_0;
wire  fifo_cout_drain_cout_drain_IO_L1_out_3_15_V_V_full_n;
assign fifo_cout_drain_cout_drain_IO_L1_out_3_15_V_V_full_n_pass_0 = fifo_cout_drain_cout_drain_IO_L1_out_3_15_V_V_full_n;
wire  cout_drain_IO_L1_out_boundary_wrapper415_U0_fifo_cout_drain_out_V_V_write;
assign cout_drain_IO_L1_out_boundary_wrapper415_U0_fifo_cout_drain_out_V_V_write = cout_drain_IO_L1_out_boundary_wrapper415_U0_fifo_cout_drain_out_V_V_write_pass_0;
wire [255:0] PE_wrapper274_U0_fifo_w_out_V_V_din;
assign PE_wrapper274_U0_fifo_w_out_V_V_din_pass_0 = PE_wrapper274_U0_fifo_w_out_V_V_din;
wire  fifo_w_PE_10_5_V_V_full_n;
reg  fifo_w_PE_10_5_V_V_full_n_q_for_broadcast;
always @ (posedge ap_clk) fifo_w_PE_10_5_V_V_full_n_q_for_broadcast <= fifo_w_PE_10_5_V_V_full_n_pass_0;
assign fifo_w_PE_10_5_V_V_full_n = fifo_w_PE_10_5_V_V_full_n_q_for_broadcast;
wire  PE_wrapper274_U0_fifo_w_out_V_V_write;
assign PE_wrapper274_U0_fifo_w_out_V_V_write_pass_0 = PE_wrapper274_U0_fifo_w_out_V_V_write;
wire [255:0] PE_wrapper262_U0_fifo_cin_out_V_V_din;
assign PE_wrapper262_U0_fifo_cin_out_V_V_din = PE_wrapper262_U0_fifo_cin_out_V_V_din_pass_1;
wire  fifo_cin_PE_10_4_V_V_full_n;
assign fifo_cin_PE_10_4_V_V_full_n_pass_1 = fifo_cin_PE_10_4_V_V_full_n;
wire  PE_wrapper262_U0_fifo_cin_out_V_V_write;
assign PE_wrapper262_U0_fifo_cin_out_V_V_write = PE_wrapper262_U0_fifo_cin_out_V_V_write_pass_1;
wire [255:0] PE_wrapper226_U0_fifo_cin_out_V_V_din;
assign PE_wrapper226_U0_fifo_cin_out_V_V_din_pass_0 = PE_wrapper226_U0_fifo_cin_out_V_V_din;
wire  fifo_cin_PE_7_4_V_V_full_n;
reg  fifo_cin_PE_7_4_V_V_full_n_q_for_broadcast;
always @ (posedge ap_clk) fifo_cin_PE_7_4_V_V_full_n_q_for_broadcast <= fifo_cin_PE_7_4_V_V_full_n_pass_0;
assign fifo_cin_PE_7_4_V_V_full_n = fifo_cin_PE_7_4_V_V_full_n_q_for_broadcast;
wire  PE_wrapper226_U0_fifo_cin_out_V_V_write;
assign PE_wrapper226_U0_fifo_cin_out_V_V_write_pass_0 = PE_wrapper226_U0_fifo_cin_out_V_V_write;
wire [31:0] PE_wrapper318_U0_fifo_cout_drain_out_V_din;
assign PE_wrapper318_U0_fifo_cout_drain_out_V_din_pass_0 = PE_wrapper318_U0_fifo_cout_drain_out_V_din;
wire  fifo_cout_drain_PE_14_0_V_full_n;
reg  fifo_cout_drain_PE_14_0_V_full_n_q_for_broadcast;
always @ (posedge ap_clk) fifo_cout_drain_PE_14_0_V_full_n_q_for_broadcast <= fifo_cout_drain_PE_14_0_V_full_n_pass_0;
assign fifo_cout_drain_PE_14_0_V_full_n = fifo_cout_drain_PE_14_0_V_full_n_q_for_broadcast;
wire  PE_wrapper318_U0_fifo_cout_drain_out_V_write;
assign PE_wrapper318_U0_fifo_cout_drain_out_V_write_pass_0 = PE_wrapper318_U0_fifo_cout_drain_out_V_write;
wire [31:0] PE_wrapper274_U0_fifo_cout_drain_out_V_din;
assign PE_wrapper274_U0_fifo_cout_drain_out_V_din_pass_0 = PE_wrapper274_U0_fifo_cout_drain_out_V_din;
wire  fifo_cout_drain_PE_10_4_V_full_n;
reg  fifo_cout_drain_PE_10_4_V_full_n_q_for_broadcast;
always @ (posedge ap_clk) fifo_cout_drain_PE_10_4_V_full_n_q_for_broadcast <= fifo_cout_drain_PE_10_4_V_full_n_pass_0;
assign fifo_cout_drain_PE_10_4_V_full_n = fifo_cout_drain_PE_10_4_V_full_n_q_for_broadcast;
wire  PE_wrapper274_U0_fifo_cout_drain_out_V_write;
assign PE_wrapper274_U0_fifo_cout_drain_out_V_write_pass_0 = PE_wrapper274_U0_fifo_cout_drain_out_V_write;
wire [31:0] PE_wrapper296_U0_fifo_cout_drain_out_V_din;
assign PE_wrapper296_U0_fifo_cout_drain_out_V_din = PE_wrapper296_U0_fifo_cout_drain_out_V_din_pass_1;
wire  fifo_cout_drain_PE_12_2_V_full_n;
assign fifo_cout_drain_PE_12_2_V_full_n_pass_1 = fifo_cout_drain_PE_12_2_V_full_n;
wire  PE_wrapper296_U0_fifo_cout_drain_out_V_write;
assign PE_wrapper296_U0_fifo_cout_drain_out_V_write = PE_wrapper296_U0_fifo_cout_drain_out_V_write_pass_1;
wire [255:0] PE_wrapper321_U0_fifo_w_out_V_V_din;
assign PE_wrapper321_U0_fifo_w_out_V_V_din_pass_0 = PE_wrapper321_U0_fifo_w_out_V_V_din;
wire  fifo_w_PE_14_4_V_V_full_n;
reg  fifo_w_PE_14_4_V_V_full_n_q_for_broadcast;
always @ (posedge ap_clk) fifo_w_PE_14_4_V_V_full_n_q_for_broadcast <= fifo_w_PE_14_4_V_V_full_n_pass_0;
assign fifo_w_PE_14_4_V_V_full_n = fifo_w_PE_14_4_V_V_full_n_q_for_broadcast;
wire  PE_wrapper321_U0_fifo_w_out_V_V_write;
assign PE_wrapper321_U0_fifo_w_out_V_V_write_pass_0 = PE_wrapper321_U0_fifo_w_out_V_V_write;
wire [31:0] PE_wrapper322_U0_fifo_cout_drain_out_V_din;
assign PE_wrapper322_U0_fifo_cout_drain_out_V_din = PE_wrapper322_U0_fifo_cout_drain_out_V_din_pass_0;
wire  fifo_cout_drain_PE_14_4_V_full_n;
assign fifo_cout_drain_PE_14_4_V_full_n_pass_0 = fifo_cout_drain_PE_14_4_V_full_n;
wire  PE_wrapper322_U0_fifo_cout_drain_out_V_write;
assign PE_wrapper322_U0_fifo_cout_drain_out_V_write = PE_wrapper322_U0_fifo_cout_drain_out_V_write_pass_0;
wire [63:0] cout_drain_IO_L1_out_wrapper401_U0_fifo_cout_drain_out_V_V_din;
assign cout_drain_IO_L1_out_wrapper401_U0_fifo_cout_drain_out_V_V_din = cout_drain_IO_L1_out_wrapper401_U0_fifo_cout_drain_out_V_V_din_pass_0;
wire  fifo_cout_drain_cout_drain_IO_L1_out_2_13_V_V_full_n;
assign fifo_cout_drain_cout_drain_IO_L1_out_2_13_V_V_full_n_pass_0 = fifo_cout_drain_cout_drain_IO_L1_out_2_13_V_V_full_n;
wire  cout_drain_IO_L1_out_wrapper401_U0_fifo_cout_drain_out_V_V_write;
assign cout_drain_IO_L1_out_wrapper401_U0_fifo_cout_drain_out_V_V_write = cout_drain_IO_L1_out_wrapper401_U0_fifo_cout_drain_out_V_V_write_pass_0;
wire [63:0] cout_drain_IO_L1_out_wrapper434_U0_fifo_cout_drain_out_V_V_din;
assign cout_drain_IO_L1_out_wrapper434_U0_fifo_cout_drain_out_V_V_din_pass_0 = cout_drain_IO_L1_out_wrapper434_U0_fifo_cout_drain_out_V_V_din;
wire  fifo_cout_drain_cout_drain_IO_L1_out_4_12_V_V_full_n;
reg  fifo_cout_drain_cout_drain_IO_L1_out_4_12_V_V_full_n_q_for_broadcast;
always @ (posedge ap_clk) fifo_cout_drain_cout_drain_IO_L1_out_4_12_V_V_full_n_q_for_broadcast <= fifo_cout_drain_cout_drain_IO_L1_out_4_12_V_V_full_n_pass_0;
assign fifo_cout_drain_cout_drain_IO_L1_out_4_12_V_V_full_n = fifo_cout_drain_cout_drain_IO_L1_out_4_12_V_V_full_n_q_for_broadcast;
wire  cout_drain_IO_L1_out_wrapper434_U0_fifo_cout_drain_out_V_V_write;
assign cout_drain_IO_L1_out_wrapper434_U0_fifo_cout_drain_out_V_V_write_pass_0 = cout_drain_IO_L1_out_wrapper434_U0_fifo_cout_drain_out_V_V_write;
wire [31:0] PE_wrapper298_U0_fifo_cout_drain_out_V_din;
assign PE_wrapper298_U0_fifo_cout_drain_out_V_din = PE_wrapper298_U0_fifo_cout_drain_out_V_din_pass_0;
wire  fifo_cout_drain_PE_12_4_V_full_n;
assign fifo_cout_drain_PE_12_4_V_full_n_pass_0 = fifo_cout_drain_PE_12_4_V_full_n;
wire  PE_wrapper298_U0_fifo_cout_drain_out_V_write;
assign PE_wrapper298_U0_fifo_cout_drain_out_V_write = PE_wrapper298_U0_fifo_cout_drain_out_V_write_pass_0;


  (* dont_touch = "yes" *) CR_X2Y6_To_CR_X3Y7 CR_X2Y6_To_CR_X3Y7_U0 (
    .PE_wrapper320_U0_fifo_cout_drain_out_V_din(PE_wrapper320_U0_fifo_cout_drain_out_V_din),
    .fifo_cout_drain_PE_14_2_V_full_n(fifo_cout_drain_PE_14_2_V_full_n),
    .PE_wrapper320_U0_fifo_cout_drain_out_V_write(PE_wrapper320_U0_fifo_cout_drain_out_V_write),
    .cout_drain_IO_L1_out_wrapper433_U0_fifo_cout_drain_out_V_V_din(cout_drain_IO_L1_out_wrapper433_U0_fifo_cout_drain_out_V_V_din),
    .fifo_cout_drain_cout_drain_IO_L1_out_4_13_V_V_full_n(fifo_cout_drain_cout_drain_IO_L1_out_4_13_V_V_full_n),
    .cout_drain_IO_L1_out_wrapper433_U0_fifo_cout_drain_out_V_V_write(cout_drain_IO_L1_out_wrapper433_U0_fifo_cout_drain_out_V_V_write),
    .PE_wrapper309_U0_fifo_cin_out_V_V_din(PE_wrapper309_U0_fifo_cin_out_V_V_din),
    .fifo_cin_PE_14_3_V_V_full_n(fifo_cin_PE_14_3_V_V_full_n),
    .PE_wrapper309_U0_fifo_cin_out_V_V_write(PE_wrapper309_U0_fifo_cin_out_V_V_write),
    .cout_drain_IO_L1_out_wrapper402_U0_fifo_cout_drain_out_V_V_din(cout_drain_IO_L1_out_wrapper402_U0_fifo_cout_drain_out_V_V_din),
    .fifo_cout_drain_cout_drain_IO_L1_out_2_12_V_V_full_n(fifo_cout_drain_cout_drain_IO_L1_out_2_12_V_V_full_n),
    .cout_drain_IO_L1_out_wrapper402_U0_fifo_cout_drain_out_V_V_write(cout_drain_IO_L1_out_wrapper402_U0_fifo_cout_drain_out_V_V_write),
    .w_IO_L2_in149_U0_fifo_w_out_V_V_din(w_IO_L2_in149_U0_fifo_w_out_V_V_din),
    .fifo_w_w_IO_L2_in_15_V_V_full_n(fifo_w_w_IO_L2_in_15_V_V_full_n),
    .w_IO_L2_in149_U0_fifo_w_out_V_V_write(w_IO_L2_in149_U0_fifo_w_out_V_V_write),
    .PE_wrapper286_U0_fifo_cout_drain_out_V_din(PE_wrapper286_U0_fifo_cout_drain_out_V_din),
    .fifo_cout_drain_PE_11_4_V_full_n(fifo_cout_drain_PE_11_4_V_full_n),
    .PE_wrapper286_U0_fifo_cout_drain_out_V_write(PE_wrapper286_U0_fifo_cout_drain_out_V_write),
    .PE_wrapper214_U0_fifo_cin_out_V_V_din(PE_wrapper214_U0_fifo_cin_out_V_V_din),
    .fifo_cin_PE_6_4_V_V_full_n(fifo_cin_PE_6_4_V_V_full_n),
    .PE_wrapper214_U0_fifo_cin_out_V_V_write(PE_wrapper214_U0_fifo_cin_out_V_V_write),
    .cout_drain_IO_L1_out_wrapper432_U0_fifo_cout_drain_out_V_V_din(cout_drain_IO_L1_out_wrapper432_U0_fifo_cout_drain_out_V_V_din),
    .fifo_cout_drain_cout_drain_IO_L1_out_4_14_V_V_full_n(fifo_cout_drain_cout_drain_IO_L1_out_4_14_V_V_full_n),
    .cout_drain_IO_L1_out_wrapper432_U0_fifo_cout_drain_out_V_V_write(cout_drain_IO_L1_out_wrapper432_U0_fifo_cout_drain_out_V_V_write),
    .PE_wrapper318_U0_fifo_w_out_V_V_din(PE_wrapper318_U0_fifo_w_out_V_V_din),
    .fifo_w_PE_14_1_V_V_full_n(fifo_w_PE_14_1_V_V_full_n),
    .PE_wrapper318_U0_fifo_w_out_V_V_write(PE_wrapper318_U0_fifo_w_out_V_V_write),
    .PE_wrapper226_U0_fifo_cout_drain_out_V_din(PE_wrapper226_U0_fifo_cout_drain_out_V_din),
    .fifo_cout_drain_PE_6_4_V_full_n(fifo_cout_drain_PE_6_4_V_full_n),
    .PE_wrapper226_U0_fifo_cout_drain_out_V_write(PE_wrapper226_U0_fifo_cout_drain_out_V_write),
    .PE_wrapper286_U0_fifo_cin_out_V_V_din(PE_wrapper286_U0_fifo_cin_out_V_V_din),
    .fifo_cin_PE_12_4_V_V_full_n(fifo_cin_PE_12_4_V_V_full_n),
    .PE_wrapper286_U0_fifo_cin_out_V_V_write(PE_wrapper286_U0_fifo_cin_out_V_V_write),
    .w_IO_L2_in148_U0_fifo_w_out_V_V_din(w_IO_L2_in148_U0_fifo_w_out_V_V_din),
    .fifo_w_w_IO_L2_in_14_V_V_full_n(fifo_w_w_IO_L2_in_14_V_V_full_n),
    .w_IO_L2_in148_U0_fifo_w_out_V_V_write(w_IO_L2_in148_U0_fifo_w_out_V_V_write),
    .PE_wrapper320_U0_fifo_cin_out_V_V_din(PE_wrapper320_U0_fifo_cin_out_V_V_din),
    .fifo_cin_PE_15_2_V_V_full_n(fifo_cin_PE_15_2_V_V_full_n),
    .PE_wrapper320_U0_fifo_cin_out_V_V_write(PE_wrapper320_U0_fifo_cin_out_V_V_write),
    .cout_drain_IO_L1_out_wrapper418_U0_fifo_cout_drain_out_V_V_din(cout_drain_IO_L1_out_wrapper418_U0_fifo_cout_drain_out_V_V_din),
    .fifo_cout_drain_cout_drain_IO_L1_out_3_12_V_V_full_n(fifo_cout_drain_cout_drain_IO_L1_out_3_12_V_V_full_n),
    .cout_drain_IO_L1_out_wrapper418_U0_fifo_cout_drain_out_V_V_write(cout_drain_IO_L1_out_wrapper418_U0_fifo_cout_drain_out_V_V_write),
    .PE_wrapper225_U0_fifo_w_out_V_V_din(PE_wrapper225_U0_fifo_w_out_V_V_din),
    .fifo_w_PE_6_4_V_V_full_n(fifo_w_PE_6_4_V_V_full_n),
    .PE_wrapper225_U0_fifo_w_out_V_V_write(PE_wrapper225_U0_fifo_w_out_V_V_write),
    .cout_drain_IO_L1_out_wrapper416_U0_fifo_cout_drain_out_V_V_din(cout_drain_IO_L1_out_wrapper416_U0_fifo_cout_drain_out_V_V_din),
    .fifo_cout_drain_cout_drain_IO_L1_out_3_14_V_V_full_n(fifo_cout_drain_cout_drain_IO_L1_out_3_14_V_V_full_n),
    .cout_drain_IO_L1_out_wrapper416_U0_fifo_cout_drain_out_V_V_write(cout_drain_IO_L1_out_wrapper416_U0_fifo_cout_drain_out_V_V_write),
    .PE_wrapper330_U0_fifo_cin_out_V_V_din(PE_wrapper330_U0_fifo_cin_out_V_V_din),
    .fifo_cin_PE_16_0_V_V_full_n(fifo_cin_PE_16_0_V_V_full_n),
    .PE_wrapper330_U0_fifo_cin_out_V_V_write(PE_wrapper330_U0_fifo_cin_out_V_V_write),
    .PE_wrapper330_U0_fifo_w_out_V_V_din(PE_wrapper330_U0_fifo_w_out_V_V_din),
    .fifo_w_PE_15_1_V_V_full_n(fifo_w_PE_15_1_V_V_full_n),
    .PE_wrapper330_U0_fifo_w_out_V_V_write(PE_wrapper330_U0_fifo_w_out_V_V_write),
    .PE_wrapper285_U0_fifo_w_out_V_V_din(PE_wrapper285_U0_fifo_w_out_V_V_din),
    .fifo_w_PE_11_4_V_V_full_n(fifo_w_PE_11_4_V_V_full_n),
    .PE_wrapper285_U0_fifo_w_out_V_V_write(PE_wrapper285_U0_fifo_w_out_V_V_write),
    .cout_drain_IO_L1_out_wrapper419_U0_fifo_cout_drain_out_V_V_din(cout_drain_IO_L1_out_wrapper419_U0_fifo_cout_drain_out_V_V_din),
    .fifo_cout_drain_cout_drain_IO_L1_out_3_11_V_V_full_n(fifo_cout_drain_cout_drain_IO_L1_out_3_11_V_V_full_n),
    .cout_drain_IO_L1_out_wrapper419_U0_fifo_cout_drain_out_V_V_write(cout_drain_IO_L1_out_wrapper419_U0_fifo_cout_drain_out_V_V_write),
    .w_IO_L2_in_boundary_U0_fifo_w_local_out_V_V_din(w_IO_L2_in_boundary_U0_fifo_w_local_out_V_V_din),
    .fifo_w_PE_15_0_V_V_full_n(fifo_w_PE_15_0_V_V_full_n),
    .w_IO_L2_in_boundary_U0_fifo_w_local_out_V_V_write(w_IO_L2_in_boundary_U0_fifo_w_local_out_V_V_write),
    .PE_wrapper273_U0_fifo_w_out_V_V_din(PE_wrapper273_U0_fifo_w_out_V_V_din),
    .fifo_w_PE_10_4_V_V_full_n(fifo_w_PE_10_4_V_V_full_n),
    .PE_wrapper273_U0_fifo_w_out_V_V_write(PE_wrapper273_U0_fifo_w_out_V_V_write),
    .PE_wrapper286_U0_fifo_w_out_V_V_din(PE_wrapper286_U0_fifo_w_out_V_V_din),
    .fifo_w_PE_11_5_V_V_full_n(fifo_w_PE_11_5_V_V_full_n),
    .PE_wrapper286_U0_fifo_w_out_V_V_write(PE_wrapper286_U0_fifo_w_out_V_V_write),
    .cout_drain_IO_L1_out_boundary_wrapper383_U0_fifo_cout_drain_out_V_V_din(cout_drain_IO_L1_out_boundary_wrapper383_U0_fifo_cout_drain_out_V_V_din),
    .fifo_cout_drain_cout_drain_IO_L1_out_1_15_V_V_full_n(fifo_cout_drain_cout_drain_IO_L1_out_1_15_V_V_full_n),
    .cout_drain_IO_L1_out_boundary_wrapper383_U0_fifo_cout_drain_out_V_V_write(cout_drain_IO_L1_out_boundary_wrapper383_U0_fifo_cout_drain_out_V_V_write),
    .PE_wrapper330_U0_fifo_cout_drain_out_V_din(PE_wrapper330_U0_fifo_cout_drain_out_V_din),
    .fifo_cout_drain_PE_15_0_V_full_n(fifo_cout_drain_PE_15_0_V_full_n),
    .PE_wrapper330_U0_fifo_cout_drain_out_V_write(PE_wrapper330_U0_fifo_cout_drain_out_V_write),
    .PE_wrapper306_U0_fifo_cin_out_V_V_din(PE_wrapper306_U0_fifo_cin_out_V_V_din),
    .fifo_cin_PE_14_0_V_V_full_n(fifo_cin_PE_14_0_V_V_full_n),
    .PE_wrapper306_U0_fifo_cin_out_V_V_write(PE_wrapper306_U0_fifo_cin_out_V_V_write),
    .PE_wrapper321_U0_fifo_cin_out_V_V_din(PE_wrapper321_U0_fifo_cin_out_V_V_din),
    .fifo_cin_PE_15_3_V_V_full_n(fifo_cin_PE_15_3_V_V_full_n),
    .PE_wrapper321_U0_fifo_cin_out_V_V_write(PE_wrapper321_U0_fifo_cin_out_V_V_write),
    .PE_wrapper285_U0_fifo_cout_drain_out_V_din(PE_wrapper285_U0_fifo_cout_drain_out_V_din),
    .fifo_cout_drain_PE_11_3_V_full_n(fifo_cout_drain_PE_11_3_V_full_n),
    .PE_wrapper285_U0_fifo_cout_drain_out_V_write(PE_wrapper285_U0_fifo_cout_drain_out_V_write),
    .PE_wrapper319_U0_fifo_w_out_V_V_din(PE_wrapper319_U0_fifo_w_out_V_V_din),
    .fifo_w_PE_14_2_V_V_full_n(fifo_w_PE_14_2_V_V_full_n),
    .PE_wrapper319_U0_fifo_w_out_V_V_write(PE_wrapper319_U0_fifo_w_out_V_V_write),
    .PE_wrapper226_U0_fifo_w_out_V_V_din(PE_wrapper226_U0_fifo_w_out_V_V_din),
    .fifo_w_PE_6_5_V_V_full_n(fifo_w_PE_6_5_V_V_full_n),
    .PE_wrapper226_U0_fifo_w_out_V_V_write(PE_wrapper226_U0_fifo_w_out_V_V_write),
    .PE_wrapper308_U0_fifo_cin_out_V_V_din(PE_wrapper308_U0_fifo_cin_out_V_V_din),
    .fifo_cin_PE_14_2_V_V_full_n(fifo_cin_PE_14_2_V_V_full_n),
    .PE_wrapper308_U0_fifo_cin_out_V_V_write(PE_wrapper308_U0_fifo_cin_out_V_V_write),
    .cout_drain_IO_L1_out_wrapper384_U0_fifo_cout_drain_out_V_V_din(cout_drain_IO_L1_out_wrapper384_U0_fifo_cout_drain_out_V_V_din),
    .fifo_cout_drain_cout_drain_IO_L1_out_1_14_V_V_full_n(fifo_cout_drain_cout_drain_IO_L1_out_1_14_V_V_full_n),
    .cout_drain_IO_L1_out_wrapper384_U0_fifo_cout_drain_out_V_V_write(cout_drain_IO_L1_out_wrapper384_U0_fifo_cout_drain_out_V_V_write),
    .PE_wrapper319_U0_fifo_cout_drain_out_V_din(PE_wrapper319_U0_fifo_cout_drain_out_V_din),
    .fifo_cout_drain_PE_14_1_V_full_n(fifo_cout_drain_PE_14_1_V_full_n),
    .PE_wrapper319_U0_fifo_cout_drain_out_V_write(PE_wrapper319_U0_fifo_cout_drain_out_V_write),
    .PE_wrapper334_U0_fifo_cout_drain_out_V_din(PE_wrapper334_U0_fifo_cout_drain_out_V_din),
    .fifo_cout_drain_PE_15_4_V_full_n(fifo_cout_drain_PE_15_4_V_full_n),
    .PE_wrapper334_U0_fifo_cout_drain_out_V_write(PE_wrapper334_U0_fifo_cout_drain_out_V_write),
    .cout_drain_IO_L1_out_boundary_wrapper415_U0_fifo_cout_drain_out_V_V_din(cout_drain_IO_L1_out_boundary_wrapper415_U0_fifo_cout_drain_out_V_V_din),
    .fifo_cout_drain_cout_drain_IO_L1_out_3_15_V_V_full_n(fifo_cout_drain_cout_drain_IO_L1_out_3_15_V_V_full_n),
    .cout_drain_IO_L1_out_boundary_wrapper415_U0_fifo_cout_drain_out_V_V_write(cout_drain_IO_L1_out_boundary_wrapper415_U0_fifo_cout_drain_out_V_V_write),
    .PE_wrapper274_U0_fifo_w_out_V_V_din(PE_wrapper274_U0_fifo_w_out_V_V_din),
    .fifo_w_PE_10_5_V_V_full_n(fifo_w_PE_10_5_V_V_full_n),
    .PE_wrapper274_U0_fifo_w_out_V_V_write(PE_wrapper274_U0_fifo_w_out_V_V_write),
    .PE_wrapper262_U0_fifo_cin_out_V_V_din(PE_wrapper262_U0_fifo_cin_out_V_V_din),
    .fifo_cin_PE_10_4_V_V_full_n(fifo_cin_PE_10_4_V_V_full_n),
    .PE_wrapper262_U0_fifo_cin_out_V_V_write(PE_wrapper262_U0_fifo_cin_out_V_V_write),
    .PE_wrapper226_U0_fifo_cin_out_V_V_din(PE_wrapper226_U0_fifo_cin_out_V_V_din),
    .fifo_cin_PE_7_4_V_V_full_n(fifo_cin_PE_7_4_V_V_full_n),
    .PE_wrapper226_U0_fifo_cin_out_V_V_write(PE_wrapper226_U0_fifo_cin_out_V_V_write),
    .PE_wrapper318_U0_fifo_cout_drain_out_V_din(PE_wrapper318_U0_fifo_cout_drain_out_V_din),
    .fifo_cout_drain_PE_14_0_V_full_n(fifo_cout_drain_PE_14_0_V_full_n),
    .PE_wrapper318_U0_fifo_cout_drain_out_V_write(PE_wrapper318_U0_fifo_cout_drain_out_V_write),
    .PE_wrapper274_U0_fifo_cout_drain_out_V_din(PE_wrapper274_U0_fifo_cout_drain_out_V_din),
    .fifo_cout_drain_PE_10_4_V_full_n(fifo_cout_drain_PE_10_4_V_full_n),
    .PE_wrapper274_U0_fifo_cout_drain_out_V_write(PE_wrapper274_U0_fifo_cout_drain_out_V_write),
    .PE_wrapper296_U0_fifo_cout_drain_out_V_din(PE_wrapper296_U0_fifo_cout_drain_out_V_din),
    .fifo_cout_drain_PE_12_2_V_full_n(fifo_cout_drain_PE_12_2_V_full_n),
    .PE_wrapper296_U0_fifo_cout_drain_out_V_write(PE_wrapper296_U0_fifo_cout_drain_out_V_write),
    .PE_wrapper321_U0_fifo_w_out_V_V_din(PE_wrapper321_U0_fifo_w_out_V_V_din),
    .fifo_w_PE_14_4_V_V_full_n(fifo_w_PE_14_4_V_V_full_n),
    .PE_wrapper321_U0_fifo_w_out_V_V_write(PE_wrapper321_U0_fifo_w_out_V_V_write),
    .PE_wrapper322_U0_fifo_cout_drain_out_V_din(PE_wrapper322_U0_fifo_cout_drain_out_V_din),
    .fifo_cout_drain_PE_14_4_V_full_n(fifo_cout_drain_PE_14_4_V_full_n),
    .PE_wrapper322_U0_fifo_cout_drain_out_V_write(PE_wrapper322_U0_fifo_cout_drain_out_V_write),
    .cout_drain_IO_L1_out_wrapper401_U0_fifo_cout_drain_out_V_V_din(cout_drain_IO_L1_out_wrapper401_U0_fifo_cout_drain_out_V_V_din),
    .fifo_cout_drain_cout_drain_IO_L1_out_2_13_V_V_full_n(fifo_cout_drain_cout_drain_IO_L1_out_2_13_V_V_full_n),
    .cout_drain_IO_L1_out_wrapper401_U0_fifo_cout_drain_out_V_V_write(cout_drain_IO_L1_out_wrapper401_U0_fifo_cout_drain_out_V_V_write),
    .cout_drain_IO_L1_out_wrapper434_U0_fifo_cout_drain_out_V_V_din(cout_drain_IO_L1_out_wrapper434_U0_fifo_cout_drain_out_V_V_din),
    .fifo_cout_drain_cout_drain_IO_L1_out_4_12_V_V_full_n(fifo_cout_drain_cout_drain_IO_L1_out_4_12_V_V_full_n),
    .cout_drain_IO_L1_out_wrapper434_U0_fifo_cout_drain_out_V_V_write(cout_drain_IO_L1_out_wrapper434_U0_fifo_cout_drain_out_V_V_write),
    .PE_wrapper298_U0_fifo_cout_drain_out_V_din(PE_wrapper298_U0_fifo_cout_drain_out_V_din),
    .fifo_cout_drain_PE_12_4_V_full_n(fifo_cout_drain_PE_12_4_V_full_n),
    .PE_wrapper298_U0_fifo_cout_drain_out_V_write(PE_wrapper298_U0_fifo_cout_drain_out_V_write),
    .ap_start(ap_start),
    .ap_done(ap_done),
    .ap_idle(ap_idle),
    .ap_ready(ap_ready),
    .ap_continue(ap_continue),
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n)
  );
endmodule


`timescale 1 ns / 1 ps
module CR_X2Y6_To_CR_X3Y7 (
  PE_wrapper320_U0_fifo_cout_drain_out_V_din,
  fifo_cout_drain_PE_14_2_V_full_n,
  PE_wrapper320_U0_fifo_cout_drain_out_V_write,
  cout_drain_IO_L1_out_wrapper433_U0_fifo_cout_drain_out_V_V_din,
  fifo_cout_drain_cout_drain_IO_L1_out_4_13_V_V_full_n,
  cout_drain_IO_L1_out_wrapper433_U0_fifo_cout_drain_out_V_V_write,
  PE_wrapper309_U0_fifo_cin_out_V_V_din,
  fifo_cin_PE_14_3_V_V_full_n,
  PE_wrapper309_U0_fifo_cin_out_V_V_write,
  cout_drain_IO_L1_out_wrapper402_U0_fifo_cout_drain_out_V_V_din,
  fifo_cout_drain_cout_drain_IO_L1_out_2_12_V_V_full_n,
  cout_drain_IO_L1_out_wrapper402_U0_fifo_cout_drain_out_V_V_write,
  w_IO_L2_in149_U0_fifo_w_out_V_V_din,
  fifo_w_w_IO_L2_in_15_V_V_full_n,
  w_IO_L2_in149_U0_fifo_w_out_V_V_write,
  PE_wrapper286_U0_fifo_cout_drain_out_V_din,
  fifo_cout_drain_PE_11_4_V_full_n,
  PE_wrapper286_U0_fifo_cout_drain_out_V_write,
  PE_wrapper214_U0_fifo_cin_out_V_V_din,
  fifo_cin_PE_6_4_V_V_full_n,
  PE_wrapper214_U0_fifo_cin_out_V_V_write,
  cout_drain_IO_L1_out_wrapper432_U0_fifo_cout_drain_out_V_V_din,
  fifo_cout_drain_cout_drain_IO_L1_out_4_14_V_V_full_n,
  cout_drain_IO_L1_out_wrapper432_U0_fifo_cout_drain_out_V_V_write,
  PE_wrapper318_U0_fifo_w_out_V_V_din,
  fifo_w_PE_14_1_V_V_full_n,
  PE_wrapper318_U0_fifo_w_out_V_V_write,
  PE_wrapper226_U0_fifo_cout_drain_out_V_din,
  fifo_cout_drain_PE_6_4_V_full_n,
  PE_wrapper226_U0_fifo_cout_drain_out_V_write,
  PE_wrapper286_U0_fifo_cin_out_V_V_din,
  fifo_cin_PE_12_4_V_V_full_n,
  PE_wrapper286_U0_fifo_cin_out_V_V_write,
  w_IO_L2_in148_U0_fifo_w_out_V_V_din,
  fifo_w_w_IO_L2_in_14_V_V_full_n,
  w_IO_L2_in148_U0_fifo_w_out_V_V_write,
  PE_wrapper320_U0_fifo_cin_out_V_V_din,
  fifo_cin_PE_15_2_V_V_full_n,
  PE_wrapper320_U0_fifo_cin_out_V_V_write,
  cout_drain_IO_L1_out_wrapper418_U0_fifo_cout_drain_out_V_V_din,
  fifo_cout_drain_cout_drain_IO_L1_out_3_12_V_V_full_n,
  cout_drain_IO_L1_out_wrapper418_U0_fifo_cout_drain_out_V_V_write,
  PE_wrapper225_U0_fifo_w_out_V_V_din,
  fifo_w_PE_6_4_V_V_full_n,
  PE_wrapper225_U0_fifo_w_out_V_V_write,
  cout_drain_IO_L1_out_wrapper416_U0_fifo_cout_drain_out_V_V_din,
  fifo_cout_drain_cout_drain_IO_L1_out_3_14_V_V_full_n,
  cout_drain_IO_L1_out_wrapper416_U0_fifo_cout_drain_out_V_V_write,
  PE_wrapper330_U0_fifo_cin_out_V_V_din,
  fifo_cin_PE_16_0_V_V_full_n,
  PE_wrapper330_U0_fifo_cin_out_V_V_write,
  PE_wrapper330_U0_fifo_w_out_V_V_din,
  fifo_w_PE_15_1_V_V_full_n,
  PE_wrapper330_U0_fifo_w_out_V_V_write,
  PE_wrapper285_U0_fifo_w_out_V_V_din,
  fifo_w_PE_11_4_V_V_full_n,
  PE_wrapper285_U0_fifo_w_out_V_V_write,
  cout_drain_IO_L1_out_wrapper419_U0_fifo_cout_drain_out_V_V_din,
  fifo_cout_drain_cout_drain_IO_L1_out_3_11_V_V_full_n,
  cout_drain_IO_L1_out_wrapper419_U0_fifo_cout_drain_out_V_V_write,
  w_IO_L2_in_boundary_U0_fifo_w_local_out_V_V_din,
  fifo_w_PE_15_0_V_V_full_n,
  w_IO_L2_in_boundary_U0_fifo_w_local_out_V_V_write,
  PE_wrapper273_U0_fifo_w_out_V_V_din,
  fifo_w_PE_10_4_V_V_full_n,
  PE_wrapper273_U0_fifo_w_out_V_V_write,
  PE_wrapper286_U0_fifo_w_out_V_V_din,
  fifo_w_PE_11_5_V_V_full_n,
  PE_wrapper286_U0_fifo_w_out_V_V_write,
  cout_drain_IO_L1_out_boundary_wrapper383_U0_fifo_cout_drain_out_V_V_din,
  fifo_cout_drain_cout_drain_IO_L1_out_1_15_V_V_full_n,
  cout_drain_IO_L1_out_boundary_wrapper383_U0_fifo_cout_drain_out_V_V_write,
  PE_wrapper330_U0_fifo_cout_drain_out_V_din,
  fifo_cout_drain_PE_15_0_V_full_n,
  PE_wrapper330_U0_fifo_cout_drain_out_V_write,
  PE_wrapper306_U0_fifo_cin_out_V_V_din,
  fifo_cin_PE_14_0_V_V_full_n,
  PE_wrapper306_U0_fifo_cin_out_V_V_write,
  PE_wrapper321_U0_fifo_cin_out_V_V_din,
  fifo_cin_PE_15_3_V_V_full_n,
  PE_wrapper321_U0_fifo_cin_out_V_V_write,
  PE_wrapper285_U0_fifo_cout_drain_out_V_din,
  fifo_cout_drain_PE_11_3_V_full_n,
  PE_wrapper285_U0_fifo_cout_drain_out_V_write,
  PE_wrapper319_U0_fifo_w_out_V_V_din,
  fifo_w_PE_14_2_V_V_full_n,
  PE_wrapper319_U0_fifo_w_out_V_V_write,
  PE_wrapper226_U0_fifo_w_out_V_V_din,
  fifo_w_PE_6_5_V_V_full_n,
  PE_wrapper226_U0_fifo_w_out_V_V_write,
  PE_wrapper308_U0_fifo_cin_out_V_V_din,
  fifo_cin_PE_14_2_V_V_full_n,
  PE_wrapper308_U0_fifo_cin_out_V_V_write,
  cout_drain_IO_L1_out_wrapper384_U0_fifo_cout_drain_out_V_V_din,
  fifo_cout_drain_cout_drain_IO_L1_out_1_14_V_V_full_n,
  cout_drain_IO_L1_out_wrapper384_U0_fifo_cout_drain_out_V_V_write,
  PE_wrapper319_U0_fifo_cout_drain_out_V_din,
  fifo_cout_drain_PE_14_1_V_full_n,
  PE_wrapper319_U0_fifo_cout_drain_out_V_write,
  PE_wrapper334_U0_fifo_cout_drain_out_V_din,
  fifo_cout_drain_PE_15_4_V_full_n,
  PE_wrapper334_U0_fifo_cout_drain_out_V_write,
  cout_drain_IO_L1_out_boundary_wrapper415_U0_fifo_cout_drain_out_V_V_din,
  fifo_cout_drain_cout_drain_IO_L1_out_3_15_V_V_full_n,
  cout_drain_IO_L1_out_boundary_wrapper415_U0_fifo_cout_drain_out_V_V_write,
  PE_wrapper274_U0_fifo_w_out_V_V_din,
  fifo_w_PE_10_5_V_V_full_n,
  PE_wrapper274_U0_fifo_w_out_V_V_write,
  PE_wrapper262_U0_fifo_cin_out_V_V_din,
  fifo_cin_PE_10_4_V_V_full_n,
  PE_wrapper262_U0_fifo_cin_out_V_V_write,
  PE_wrapper226_U0_fifo_cin_out_V_V_din,
  fifo_cin_PE_7_4_V_V_full_n,
  PE_wrapper226_U0_fifo_cin_out_V_V_write,
  PE_wrapper318_U0_fifo_cout_drain_out_V_din,
  fifo_cout_drain_PE_14_0_V_full_n,
  PE_wrapper318_U0_fifo_cout_drain_out_V_write,
  PE_wrapper274_U0_fifo_cout_drain_out_V_din,
  fifo_cout_drain_PE_10_4_V_full_n,
  PE_wrapper274_U0_fifo_cout_drain_out_V_write,
  PE_wrapper296_U0_fifo_cout_drain_out_V_din,
  fifo_cout_drain_PE_12_2_V_full_n,
  PE_wrapper296_U0_fifo_cout_drain_out_V_write,
  PE_wrapper321_U0_fifo_w_out_V_V_din,
  fifo_w_PE_14_4_V_V_full_n,
  PE_wrapper321_U0_fifo_w_out_V_V_write,
  PE_wrapper322_U0_fifo_cout_drain_out_V_din,
  fifo_cout_drain_PE_14_4_V_full_n,
  PE_wrapper322_U0_fifo_cout_drain_out_V_write,
  cout_drain_IO_L1_out_wrapper401_U0_fifo_cout_drain_out_V_V_din,
  fifo_cout_drain_cout_drain_IO_L1_out_2_13_V_V_full_n,
  cout_drain_IO_L1_out_wrapper401_U0_fifo_cout_drain_out_V_V_write,
  cout_drain_IO_L1_out_wrapper434_U0_fifo_cout_drain_out_V_V_din,
  fifo_cout_drain_cout_drain_IO_L1_out_4_12_V_V_full_n,
  cout_drain_IO_L1_out_wrapper434_U0_fifo_cout_drain_out_V_V_write,
  PE_wrapper298_U0_fifo_cout_drain_out_V_din,
  fifo_cout_drain_PE_12_4_V_full_n,
  PE_wrapper298_U0_fifo_cout_drain_out_V_write,
  ap_start,
  ap_done,
  ap_idle,
  ap_ready,
  ap_continue,
  ap_clk,
  ap_rst_n
);
parameter C_S_AXI_CONTROL_DATA_WIDTH = 32;
parameter C_S_AXI_CONTROL_ADDR_WIDTH = 6;
parameter C_S_AXI_DATA_WIDTH = 32;
parameter C_S_AXI_ADDR_WIDTH = 32;
parameter C_M_AXI_GMEM_CIN_ID_WIDTH = 1;
parameter C_M_AXI_GMEM_CIN_ADDR_WIDTH = 64;
parameter C_M_AXI_GMEM_CIN_DATA_WIDTH = 512;
parameter C_M_AXI_GMEM_CIN_AWUSER_WIDTH = 1;
parameter C_M_AXI_GMEM_CIN_ARUSER_WIDTH = 1;
parameter C_M_AXI_GMEM_CIN_WUSER_WIDTH = 1;
parameter C_M_AXI_GMEM_CIN_RUSER_WIDTH = 1;
parameter C_M_AXI_GMEM_CIN_BUSER_WIDTH = 1;
parameter C_M_AXI_GMEM_CIN_USER_VALUE = 0;
parameter C_M_AXI_GMEM_CIN_PROT_VALUE = 0;
parameter C_M_AXI_GMEM_CIN_CACHE_VALUE = 3;
parameter C_M_AXI_ID_WIDTH = 1;
parameter C_M_AXI_ADDR_WIDTH = 64;
parameter C_M_AXI_DATA_WIDTH = 32;
parameter C_M_AXI_AWUSER_WIDTH = 1;
parameter C_M_AXI_ARUSER_WIDTH = 1;
parameter C_M_AXI_WUSER_WIDTH = 1;
parameter C_M_AXI_RUSER_WIDTH = 1;
parameter C_M_AXI_BUSER_WIDTH = 1;
parameter C_M_AXI_GMEM_COUT_ID_WIDTH = 1;
parameter C_M_AXI_GMEM_COUT_ADDR_WIDTH = 64;
parameter C_M_AXI_GMEM_COUT_DATA_WIDTH = 512;
parameter C_M_AXI_GMEM_COUT_AWUSER_WIDTH = 1;
parameter C_M_AXI_GMEM_COUT_ARUSER_WIDTH = 1;
parameter C_M_AXI_GMEM_COUT_WUSER_WIDTH = 1;
parameter C_M_AXI_GMEM_COUT_RUSER_WIDTH = 1;
parameter C_M_AXI_GMEM_COUT_BUSER_WIDTH = 1;
parameter C_M_AXI_GMEM_COUT_USER_VALUE = 0;
parameter C_M_AXI_GMEM_COUT_PROT_VALUE = 0;
parameter C_M_AXI_GMEM_COUT_CACHE_VALUE = 3;
parameter C_M_AXI_GMEM_W_ID_WIDTH = 1;
parameter C_M_AXI_GMEM_W_ADDR_WIDTH = 64;
parameter C_M_AXI_GMEM_W_DATA_WIDTH = 512;
parameter C_M_AXI_GMEM_W_AWUSER_WIDTH = 1;
parameter C_M_AXI_GMEM_W_ARUSER_WIDTH = 1;
parameter C_M_AXI_GMEM_W_WUSER_WIDTH = 1;
parameter C_M_AXI_GMEM_W_RUSER_WIDTH = 1;
parameter C_M_AXI_GMEM_W_BUSER_WIDTH = 1;
parameter C_M_AXI_GMEM_W_USER_VALUE = 0;
parameter C_M_AXI_GMEM_W_PROT_VALUE = 0;
parameter C_M_AXI_GMEM_W_CACHE_VALUE = 3;
parameter C_S_AXI_CONTROL_WSTRB_WIDTH = 32 / 8;
parameter C_S_AXI_WSTRB_WIDTH = 32 / 8;
parameter C_M_AXI_GMEM_CIN_WSTRB_WIDTH = 512 / 8;
parameter C_M_AXI_WSTRB_WIDTH = 32 / 8;
parameter C_M_AXI_GMEM_COUT_WSTRB_WIDTH = 512 / 8;
parameter C_M_AXI_GMEM_W_WSTRB_WIDTH = 512 / 8;
reg ap_rst_n_inv;
wire w_IO_L2_in149_U0_ap_start;
wire w_IO_L2_in149_U0_ap_done;
wire w_IO_L2_in149_U0_ap_continue;
wire w_IO_L2_in149_U0_ap_idle;
wire w_IO_L2_in149_U0_ap_ready;
wire w_IO_L2_in149_U0_fifo_w_in_V_V_read;
wire [255:0] w_IO_L2_in149_U0_fifo_w_local_out_V_V_din;
wire w_IO_L2_in149_U0_fifo_w_local_out_V_V_write;
wire PE_wrapper226_U0_ap_start;
wire PE_wrapper226_U0_ap_done;
wire PE_wrapper226_U0_ap_continue;
wire PE_wrapper226_U0_ap_idle;
wire PE_wrapper226_U0_ap_ready;
wire PE_wrapper226_U0_fifo_cin_in_V_V_read;
wire PE_wrapper226_U0_fifo_w_in_V_V_read;
wire PE_wrapper274_U0_ap_start;
wire PE_wrapper274_U0_ap_done;
wire PE_wrapper274_U0_ap_continue;
wire PE_wrapper274_U0_ap_idle;
wire PE_wrapper274_U0_ap_ready;
wire PE_wrapper274_U0_fifo_cin_in_V_V_read;
wire [255:0] PE_wrapper274_U0_fifo_cin_out_V_V_din;
wire PE_wrapper274_U0_fifo_cin_out_V_V_write;
wire PE_wrapper274_U0_fifo_w_in_V_V_read;
wire PE_wrapper286_U0_ap_start;
wire PE_wrapper286_U0_ap_done;
wire PE_wrapper286_U0_ap_continue;
wire PE_wrapper286_U0_ap_idle;
wire PE_wrapper286_U0_ap_ready;
wire PE_wrapper286_U0_fifo_cin_in_V_V_read;
wire PE_wrapper286_U0_fifo_w_in_V_V_read;
wire PE_wrapper318_U0_ap_start;
wire PE_wrapper318_U0_ap_done;
wire PE_wrapper318_U0_ap_continue;
wire PE_wrapper318_U0_ap_idle;
wire PE_wrapper318_U0_ap_ready;
wire PE_wrapper318_U0_fifo_cin_in_V_V_read;
wire [255:0] PE_wrapper318_U0_fifo_cin_out_V_V_din;
wire PE_wrapper318_U0_fifo_cin_out_V_V_write;
wire PE_wrapper318_U0_fifo_w_in_V_V_read;
wire PE_wrapper320_U0_ap_start;
wire PE_wrapper320_U0_ap_done;
wire PE_wrapper320_U0_ap_continue;
wire PE_wrapper320_U0_ap_idle;
wire PE_wrapper320_U0_ap_ready;
wire PE_wrapper320_U0_fifo_cin_in_V_V_read;
wire PE_wrapper320_U0_fifo_w_in_V_V_read;
wire [255:0] PE_wrapper320_U0_fifo_w_out_V_V_din;
wire PE_wrapper320_U0_fifo_w_out_V_V_write;
wire PE_wrapper321_U0_ap_start;
wire PE_wrapper321_U0_ap_done;
wire PE_wrapper321_U0_ap_continue;
wire PE_wrapper321_U0_ap_idle;
wire PE_wrapper321_U0_ap_ready;
wire PE_wrapper321_U0_fifo_cin_in_V_V_read;
wire [31:0] PE_wrapper321_U0_fifo_cout_drain_out_V_din;
wire PE_wrapper321_U0_fifo_cout_drain_out_V_write;
wire PE_wrapper321_U0_fifo_w_in_V_V_read;
wire PE_wrapper330_U0_ap_start;
wire PE_wrapper330_U0_ap_done;
wire PE_wrapper330_U0_ap_continue;
wire PE_wrapper330_U0_ap_idle;
wire PE_wrapper330_U0_ap_ready;
wire PE_wrapper330_U0_fifo_cin_in_V_V_read;
wire PE_wrapper330_U0_fifo_w_in_V_V_read;
wire cout_drain_IO_L1_out_wrapper384_U0_ap_start;
wire cout_drain_IO_L1_out_wrapper384_U0_ap_done;
wire cout_drain_IO_L1_out_wrapper384_U0_ap_continue;
wire cout_drain_IO_L1_out_wrapper384_U0_ap_idle;
wire cout_drain_IO_L1_out_wrapper384_U0_ap_ready;
wire cout_drain_IO_L1_out_wrapper384_U0_fifo_cout_drain_in_V_V_read;
wire cout_drain_IO_L1_out_wrapper384_U0_fifo_cout_drain_local_in_V_read;
wire cout_drain_IO_L1_out_wrapper402_U0_ap_start;
wire cout_drain_IO_L1_out_wrapper402_U0_ap_done;
wire cout_drain_IO_L1_out_wrapper402_U0_ap_continue;
wire cout_drain_IO_L1_out_wrapper402_U0_ap_idle;
wire cout_drain_IO_L1_out_wrapper402_U0_ap_ready;
wire cout_drain_IO_L1_out_wrapper402_U0_fifo_cout_drain_in_V_V_read;
wire cout_drain_IO_L1_out_wrapper402_U0_fifo_cout_drain_local_in_V_read;
wire cout_drain_IO_L1_out_wrapper416_U0_ap_start;
wire cout_drain_IO_L1_out_wrapper416_U0_ap_done;
wire cout_drain_IO_L1_out_wrapper416_U0_ap_continue;
wire cout_drain_IO_L1_out_wrapper416_U0_ap_idle;
wire cout_drain_IO_L1_out_wrapper416_U0_ap_ready;
wire cout_drain_IO_L1_out_wrapper416_U0_fifo_cout_drain_in_V_V_read;
wire cout_drain_IO_L1_out_wrapper416_U0_fifo_cout_drain_local_in_V_read;
wire cout_drain_IO_L1_out_wrapper419_U0_ap_start;
wire cout_drain_IO_L1_out_wrapper419_U0_ap_done;
wire cout_drain_IO_L1_out_wrapper419_U0_ap_continue;
wire cout_drain_IO_L1_out_wrapper419_U0_ap_idle;
wire cout_drain_IO_L1_out_wrapper419_U0_ap_ready;
wire cout_drain_IO_L1_out_wrapper419_U0_fifo_cout_drain_in_V_V_read;
wire cout_drain_IO_L1_out_wrapper419_U0_fifo_cout_drain_local_in_V_read;
wire cout_drain_IO_L1_out_boundary_wrapper431_U0_ap_start;
wire cout_drain_IO_L1_out_boundary_wrapper431_U0_ap_done;
wire cout_drain_IO_L1_out_boundary_wrapper431_U0_ap_continue;
wire cout_drain_IO_L1_out_boundary_wrapper431_U0_ap_idle;
wire cout_drain_IO_L1_out_boundary_wrapper431_U0_ap_ready;
wire [63:0] cout_drain_IO_L1_out_boundary_wrapper431_U0_fifo_cout_drain_out_V_V_din;
wire cout_drain_IO_L1_out_boundary_wrapper431_U0_fifo_cout_drain_out_V_V_write;
wire cout_drain_IO_L1_out_boundary_wrapper431_U0_fifo_cout_drain_local_in_V_read;
wire cout_drain_IO_L1_out_wrapper432_U0_ap_start;
wire cout_drain_IO_L1_out_wrapper432_U0_ap_done;
wire cout_drain_IO_L1_out_wrapper432_U0_ap_continue;
wire cout_drain_IO_L1_out_wrapper432_U0_ap_idle;
wire cout_drain_IO_L1_out_wrapper432_U0_ap_ready;
wire cout_drain_IO_L1_out_wrapper432_U0_fifo_cout_drain_in_V_V_read;
wire cout_drain_IO_L1_out_wrapper432_U0_fifo_cout_drain_local_in_V_read;
wire cout_drain_IO_L1_out_wrapper434_U0_ap_start;
wire cout_drain_IO_L1_out_wrapper434_U0_ap_done;
wire cout_drain_IO_L1_out_wrapper434_U0_ap_continue;
wire cout_drain_IO_L1_out_wrapper434_U0_ap_idle;
wire cout_drain_IO_L1_out_wrapper434_U0_ap_ready;
wire cout_drain_IO_L1_out_wrapper434_U0_fifo_cout_drain_in_V_V_read;
wire cout_drain_IO_L1_out_wrapper434_U0_fifo_cout_drain_local_in_V_read;
wire [255:0] fifo_w_w_IO_L2_in_14_V_V_dout;
wire fifo_w_w_IO_L2_in_14_V_V_empty_n;
wire fifo_w_PE_14_0_V_V_full_n;
wire [255:0] fifo_w_PE_14_0_V_V_dout;
wire fifo_w_PE_14_0_V_V_empty_n;
wire [255:0] fifo_w_PE_15_0_V_V_dout;
wire fifo_w_PE_15_0_V_V_empty_n;
wire [255:0] fifo_cin_PE_6_4_V_V_dout;
wire fifo_cin_PE_6_4_V_V_empty_n;
wire [255:0] fifo_w_PE_6_4_V_V_dout;
wire fifo_w_PE_6_4_V_V_empty_n;
wire [255:0] fifo_cin_PE_10_4_V_V_dout;
wire fifo_cin_PE_10_4_V_V_empty_n;
wire [255:0] fifo_w_PE_10_4_V_V_dout;
wire fifo_w_PE_10_4_V_V_empty_n;
wire fifo_cin_PE_11_4_V_V_full_n;
wire [255:0] fifo_cin_PE_11_4_V_V_dout;
wire fifo_cin_PE_11_4_V_V_empty_n;
wire [31:0] fifo_cout_drain_PE_11_3_V_dout;
wire fifo_cout_drain_PE_11_3_V_empty_n;
wire [255:0] fifo_w_PE_11_4_V_V_dout;
wire fifo_w_PE_11_4_V_V_empty_n;
wire [31:0] fifo_cout_drain_PE_12_2_V_dout;
wire fifo_cout_drain_PE_12_2_V_empty_n;
wire [31:0] fifo_cout_drain_PE_12_4_V_dout;
wire fifo_cout_drain_PE_12_4_V_empty_n;
wire [255:0] fifo_cin_PE_14_0_V_V_dout;
wire fifo_cin_PE_14_0_V_V_empty_n;
wire [255:0] fifo_cin_PE_14_2_V_V_dout;
wire fifo_cin_PE_14_2_V_V_empty_n;
wire [255:0] fifo_cin_PE_14_3_V_V_dout;
wire fifo_cin_PE_14_3_V_V_empty_n;
wire fifo_cin_PE_15_0_V_V_full_n;
wire [255:0] fifo_cin_PE_15_0_V_V_dout;
wire fifo_cin_PE_15_0_V_V_empty_n;
wire [31:0] fifo_cout_drain_PE_14_1_V_dout;
wire fifo_cout_drain_PE_14_1_V_empty_n;
wire [255:0] fifo_w_PE_14_2_V_V_dout;
wire fifo_w_PE_14_2_V_V_empty_n;
wire fifo_w_PE_14_3_V_V_full_n;
wire [255:0] fifo_w_PE_14_3_V_V_dout;
wire fifo_w_PE_14_3_V_V_empty_n;
wire fifo_cout_drain_PE_14_3_V_full_n;
wire [31:0] fifo_cout_drain_PE_14_3_V_dout;
wire fifo_cout_drain_PE_14_3_V_empty_n;
wire [31:0] fifo_cout_drain_PE_14_4_V_dout;
wire fifo_cout_drain_PE_14_4_V_empty_n;
wire [31:0] fifo_cout_drain_PE_15_4_V_dout;
wire fifo_cout_drain_PE_15_4_V_empty_n;
wire [63:0] fifo_cout_drain_cout_drain_IO_L1_out_1_15_V_V_dout;
wire fifo_cout_drain_cout_drain_IO_L1_out_1_15_V_V_empty_n;
wire [63:0] fifo_cout_drain_cout_drain_IO_L1_out_2_13_V_V_dout;
wire fifo_cout_drain_cout_drain_IO_L1_out_2_13_V_V_empty_n;
wire [63:0] fifo_cout_drain_cout_drain_IO_L1_out_3_15_V_V_dout;
wire fifo_cout_drain_cout_drain_IO_L1_out_3_15_V_V_empty_n;
wire [63:0] fifo_cout_drain_cout_drain_IO_L1_out_3_12_V_V_dout;
wire fifo_cout_drain_cout_drain_IO_L1_out_3_12_V_V_empty_n;
wire fifo_cout_drain_cout_drain_IO_L1_out_4_15_V_V_full_n;
wire [63:0] fifo_cout_drain_cout_drain_IO_L1_out_4_15_V_V_dout;
wire fifo_cout_drain_cout_drain_IO_L1_out_4_15_V_V_empty_n;
wire [63:0] fifo_cout_drain_cout_drain_IO_L1_out_4_13_V_V_dout;
wire fifo_cout_drain_cout_drain_IO_L1_out_4_13_V_V_empty_n;
// pipeline ap_start
(* shreg_extract = "no" *) reg ap_start_p1;
(* shreg_extract = "no" *) reg ap_start_p2;
(* shreg_extract = "no" *) reg ap_start_pipe;
// pipeline ap_rst_n
(* shreg_extract = "no" *) reg ap_rst_p1;
(* shreg_extract = "no" *) reg ap_rst_p2;
(* shreg_extract = "no" *) reg ap_rst_pipe;
(* shreg_extract = "no" *) reg ap_rst_n_p1;
(* shreg_extract = "no" *) reg ap_rst_n_p2;
(* shreg_extract = "no" *) reg ap_rst_n_pipe;
output [31:0] PE_wrapper320_U0_fifo_cout_drain_out_V_din;
input  fifo_cout_drain_PE_14_2_V_full_n;
output  PE_wrapper320_U0_fifo_cout_drain_out_V_write;
input [63:0] cout_drain_IO_L1_out_wrapper433_U0_fifo_cout_drain_out_V_V_din;
output  fifo_cout_drain_cout_drain_IO_L1_out_4_13_V_V_full_n;
input  cout_drain_IO_L1_out_wrapper433_U0_fifo_cout_drain_out_V_V_write;
input [255:0] PE_wrapper309_U0_fifo_cin_out_V_V_din;
output  fifo_cin_PE_14_3_V_V_full_n;
input  PE_wrapper309_U0_fifo_cin_out_V_V_write;
output [63:0] cout_drain_IO_L1_out_wrapper402_U0_fifo_cout_drain_out_V_V_din;
input  fifo_cout_drain_cout_drain_IO_L1_out_2_12_V_V_full_n;
output  cout_drain_IO_L1_out_wrapper402_U0_fifo_cout_drain_out_V_V_write;
output [255:0] w_IO_L2_in149_U0_fifo_w_out_V_V_din;
input  fifo_w_w_IO_L2_in_15_V_V_full_n;
output  w_IO_L2_in149_U0_fifo_w_out_V_V_write;
output [31:0] PE_wrapper286_U0_fifo_cout_drain_out_V_din;
input  fifo_cout_drain_PE_11_4_V_full_n;
output  PE_wrapper286_U0_fifo_cout_drain_out_V_write;
input [255:0] PE_wrapper214_U0_fifo_cin_out_V_V_din;
output  fifo_cin_PE_6_4_V_V_full_n;
input  PE_wrapper214_U0_fifo_cin_out_V_V_write;
output [63:0] cout_drain_IO_L1_out_wrapper432_U0_fifo_cout_drain_out_V_V_din;
input  fifo_cout_drain_cout_drain_IO_L1_out_4_14_V_V_full_n;
output  cout_drain_IO_L1_out_wrapper432_U0_fifo_cout_drain_out_V_V_write;
output [255:0] PE_wrapper318_U0_fifo_w_out_V_V_din;
input  fifo_w_PE_14_1_V_V_full_n;
output  PE_wrapper318_U0_fifo_w_out_V_V_write;
output [31:0] PE_wrapper226_U0_fifo_cout_drain_out_V_din;
input  fifo_cout_drain_PE_6_4_V_full_n;
output  PE_wrapper226_U0_fifo_cout_drain_out_V_write;
output [255:0] PE_wrapper286_U0_fifo_cin_out_V_V_din;
input  fifo_cin_PE_12_4_V_V_full_n;
output  PE_wrapper286_U0_fifo_cin_out_V_V_write;
input [255:0] w_IO_L2_in148_U0_fifo_w_out_V_V_din;
output  fifo_w_w_IO_L2_in_14_V_V_full_n;
input  w_IO_L2_in148_U0_fifo_w_out_V_V_write;
output [255:0] PE_wrapper320_U0_fifo_cin_out_V_V_din;
input  fifo_cin_PE_15_2_V_V_full_n;
output  PE_wrapper320_U0_fifo_cin_out_V_V_write;
input [63:0] cout_drain_IO_L1_out_wrapper418_U0_fifo_cout_drain_out_V_V_din;
output  fifo_cout_drain_cout_drain_IO_L1_out_3_12_V_V_full_n;
input  cout_drain_IO_L1_out_wrapper418_U0_fifo_cout_drain_out_V_V_write;
input [255:0] PE_wrapper225_U0_fifo_w_out_V_V_din;
output  fifo_w_PE_6_4_V_V_full_n;
input  PE_wrapper225_U0_fifo_w_out_V_V_write;
output [63:0] cout_drain_IO_L1_out_wrapper416_U0_fifo_cout_drain_out_V_V_din;
input  fifo_cout_drain_cout_drain_IO_L1_out_3_14_V_V_full_n;
output  cout_drain_IO_L1_out_wrapper416_U0_fifo_cout_drain_out_V_V_write;
output [255:0] PE_wrapper330_U0_fifo_cin_out_V_V_din;
input  fifo_cin_PE_16_0_V_V_full_n;
output  PE_wrapper330_U0_fifo_cin_out_V_V_write;
output [255:0] PE_wrapper330_U0_fifo_w_out_V_V_din;
input  fifo_w_PE_15_1_V_V_full_n;
output  PE_wrapper330_U0_fifo_w_out_V_V_write;
input [255:0] PE_wrapper285_U0_fifo_w_out_V_V_din;
output  fifo_w_PE_11_4_V_V_full_n;
input  PE_wrapper285_U0_fifo_w_out_V_V_write;
output [63:0] cout_drain_IO_L1_out_wrapper419_U0_fifo_cout_drain_out_V_V_din;
input  fifo_cout_drain_cout_drain_IO_L1_out_3_11_V_V_full_n;
output  cout_drain_IO_L1_out_wrapper419_U0_fifo_cout_drain_out_V_V_write;
input [255:0] w_IO_L2_in_boundary_U0_fifo_w_local_out_V_V_din;
output  fifo_w_PE_15_0_V_V_full_n;
input  w_IO_L2_in_boundary_U0_fifo_w_local_out_V_V_write;
input [255:0] PE_wrapper273_U0_fifo_w_out_V_V_din;
output  fifo_w_PE_10_4_V_V_full_n;
input  PE_wrapper273_U0_fifo_w_out_V_V_write;
output [255:0] PE_wrapper286_U0_fifo_w_out_V_V_din;
input  fifo_w_PE_11_5_V_V_full_n;
output  PE_wrapper286_U0_fifo_w_out_V_V_write;
input [63:0] cout_drain_IO_L1_out_boundary_wrapper383_U0_fifo_cout_drain_out_V_V_din;
output  fifo_cout_drain_cout_drain_IO_L1_out_1_15_V_V_full_n;
input  cout_drain_IO_L1_out_boundary_wrapper383_U0_fifo_cout_drain_out_V_V_write;
output [31:0] PE_wrapper330_U0_fifo_cout_drain_out_V_din;
input  fifo_cout_drain_PE_15_0_V_full_n;
output  PE_wrapper330_U0_fifo_cout_drain_out_V_write;
input [255:0] PE_wrapper306_U0_fifo_cin_out_V_V_din;
output  fifo_cin_PE_14_0_V_V_full_n;
input  PE_wrapper306_U0_fifo_cin_out_V_V_write;
output [255:0] PE_wrapper321_U0_fifo_cin_out_V_V_din;
input  fifo_cin_PE_15_3_V_V_full_n;
output  PE_wrapper321_U0_fifo_cin_out_V_V_write;
input [31:0] PE_wrapper285_U0_fifo_cout_drain_out_V_din;
output  fifo_cout_drain_PE_11_3_V_full_n;
input  PE_wrapper285_U0_fifo_cout_drain_out_V_write;
input [255:0] PE_wrapper319_U0_fifo_w_out_V_V_din;
output  fifo_w_PE_14_2_V_V_full_n;
input  PE_wrapper319_U0_fifo_w_out_V_V_write;
output [255:0] PE_wrapper226_U0_fifo_w_out_V_V_din;
input  fifo_w_PE_6_5_V_V_full_n;
output  PE_wrapper226_U0_fifo_w_out_V_V_write;
input [255:0] PE_wrapper308_U0_fifo_cin_out_V_V_din;
output  fifo_cin_PE_14_2_V_V_full_n;
input  PE_wrapper308_U0_fifo_cin_out_V_V_write;
output [63:0] cout_drain_IO_L1_out_wrapper384_U0_fifo_cout_drain_out_V_V_din;
input  fifo_cout_drain_cout_drain_IO_L1_out_1_14_V_V_full_n;
output  cout_drain_IO_L1_out_wrapper384_U0_fifo_cout_drain_out_V_V_write;
input [31:0] PE_wrapper319_U0_fifo_cout_drain_out_V_din;
output  fifo_cout_drain_PE_14_1_V_full_n;
input  PE_wrapper319_U0_fifo_cout_drain_out_V_write;
input [31:0] PE_wrapper334_U0_fifo_cout_drain_out_V_din;
output  fifo_cout_drain_PE_15_4_V_full_n;
input  PE_wrapper334_U0_fifo_cout_drain_out_V_write;
input [63:0] cout_drain_IO_L1_out_boundary_wrapper415_U0_fifo_cout_drain_out_V_V_din;
output  fifo_cout_drain_cout_drain_IO_L1_out_3_15_V_V_full_n;
input  cout_drain_IO_L1_out_boundary_wrapper415_U0_fifo_cout_drain_out_V_V_write;
output [255:0] PE_wrapper274_U0_fifo_w_out_V_V_din;
input  fifo_w_PE_10_5_V_V_full_n;
output  PE_wrapper274_U0_fifo_w_out_V_V_write;
input [255:0] PE_wrapper262_U0_fifo_cin_out_V_V_din;
output  fifo_cin_PE_10_4_V_V_full_n;
input  PE_wrapper262_U0_fifo_cin_out_V_V_write;
output [255:0] PE_wrapper226_U0_fifo_cin_out_V_V_din;
input  fifo_cin_PE_7_4_V_V_full_n;
output  PE_wrapper226_U0_fifo_cin_out_V_V_write;
output [31:0] PE_wrapper318_U0_fifo_cout_drain_out_V_din;
input  fifo_cout_drain_PE_14_0_V_full_n;
output  PE_wrapper318_U0_fifo_cout_drain_out_V_write;
output [31:0] PE_wrapper274_U0_fifo_cout_drain_out_V_din;
input  fifo_cout_drain_PE_10_4_V_full_n;
output  PE_wrapper274_U0_fifo_cout_drain_out_V_write;
input [31:0] PE_wrapper296_U0_fifo_cout_drain_out_V_din;
output  fifo_cout_drain_PE_12_2_V_full_n;
input  PE_wrapper296_U0_fifo_cout_drain_out_V_write;
output [255:0] PE_wrapper321_U0_fifo_w_out_V_V_din;
input  fifo_w_PE_14_4_V_V_full_n;
output  PE_wrapper321_U0_fifo_w_out_V_V_write;
input [31:0] PE_wrapper322_U0_fifo_cout_drain_out_V_din;
output  fifo_cout_drain_PE_14_4_V_full_n;
input  PE_wrapper322_U0_fifo_cout_drain_out_V_write;
input [63:0] cout_drain_IO_L1_out_wrapper401_U0_fifo_cout_drain_out_V_V_din;
output  fifo_cout_drain_cout_drain_IO_L1_out_2_13_V_V_full_n;
input  cout_drain_IO_L1_out_wrapper401_U0_fifo_cout_drain_out_V_V_write;
output [63:0] cout_drain_IO_L1_out_wrapper434_U0_fifo_cout_drain_out_V_V_din;
input  fifo_cout_drain_cout_drain_IO_L1_out_4_12_V_V_full_n;
output  cout_drain_IO_L1_out_wrapper434_U0_fifo_cout_drain_out_V_V_write;
input [31:0] PE_wrapper298_U0_fifo_cout_drain_out_V_din;
output  fifo_cout_drain_PE_12_4_V_full_n;
input  PE_wrapper298_U0_fifo_cout_drain_out_V_write;
input  ap_start;
output ap_done;
output ap_idle;
output ap_ready;
input  ap_continue;
input ap_clk;
input ap_rst_n;
(* keep_hierarchy = "yes" *)
kernel0_w_IO_L2_in149
w_IO_L2_in149_U0
(
  .ap_clk(ap_clk),
  .ap_rst(ap_rst_pipe),
  .ap_start(ap_start_pipe),
  .ap_done(w_IO_L2_in149_U0_ap_done),
  .ap_continue(1'b1),
  .ap_idle(w_IO_L2_in149_U0_ap_idle),
  .ap_ready(w_IO_L2_in149_U0_ap_ready),
  .fifo_w_in_V_V_dout(fifo_w_w_IO_L2_in_14_V_V_dout),
  .fifo_w_in_V_V_empty_n(fifo_w_w_IO_L2_in_14_V_V_empty_n),
  .fifo_w_in_V_V_read(w_IO_L2_in149_U0_fifo_w_in_V_V_read),
  .fifo_w_out_V_V_din(w_IO_L2_in149_U0_fifo_w_out_V_V_din),
  .fifo_w_out_V_V_full_n(fifo_w_w_IO_L2_in_15_V_V_full_n),
  .fifo_w_out_V_V_write(w_IO_L2_in149_U0_fifo_w_out_V_V_write),
  .fifo_w_local_out_V_V_din(w_IO_L2_in149_U0_fifo_w_local_out_V_V_din),
  .fifo_w_local_out_V_V_full_n(fifo_w_PE_14_0_V_V_full_n),
  .fifo_w_local_out_V_V_write(w_IO_L2_in149_U0_fifo_w_local_out_V_V_write)
);

(* keep_hierarchy = "yes" *)
kernel0_PE_wrapper226
PE_wrapper226_U0
(
  .ap_clk(ap_clk),
  .ap_rst(ap_rst_pipe),
  .ap_start(ap_start_pipe),
  .ap_done(PE_wrapper226_U0_ap_done),
  .ap_continue(1'b1),
  .ap_idle(PE_wrapper226_U0_ap_idle),
  .ap_ready(PE_wrapper226_U0_ap_ready),
  .fifo_cin_in_V_V_dout(fifo_cin_PE_6_4_V_V_dout),
  .fifo_cin_in_V_V_empty_n(fifo_cin_PE_6_4_V_V_empty_n),
  .fifo_cin_in_V_V_read(PE_wrapper226_U0_fifo_cin_in_V_V_read),
  .fifo_cin_out_V_V_din(PE_wrapper226_U0_fifo_cin_out_V_V_din),
  .fifo_cin_out_V_V_full_n(fifo_cin_PE_7_4_V_V_full_n),
  .fifo_cin_out_V_V_write(PE_wrapper226_U0_fifo_cin_out_V_V_write),
  .fifo_cout_drain_out_V_din(PE_wrapper226_U0_fifo_cout_drain_out_V_din),
  .fifo_cout_drain_out_V_full_n(fifo_cout_drain_PE_6_4_V_full_n),
  .fifo_cout_drain_out_V_write(PE_wrapper226_U0_fifo_cout_drain_out_V_write),
  .fifo_w_in_V_V_dout(fifo_w_PE_6_4_V_V_dout),
  .fifo_w_in_V_V_empty_n(fifo_w_PE_6_4_V_V_empty_n),
  .fifo_w_in_V_V_read(PE_wrapper226_U0_fifo_w_in_V_V_read),
  .fifo_w_out_V_V_din(PE_wrapper226_U0_fifo_w_out_V_V_din),
  .fifo_w_out_V_V_full_n(fifo_w_PE_6_5_V_V_full_n),
  .fifo_w_out_V_V_write(PE_wrapper226_U0_fifo_w_out_V_V_write)
);

(* keep_hierarchy = "yes" *)
kernel0_PE_wrapper274
PE_wrapper274_U0
(
  .ap_clk(ap_clk),
  .ap_rst(ap_rst_pipe),
  .ap_start(ap_start_pipe),
  .ap_done(PE_wrapper274_U0_ap_done),
  .ap_continue(1'b1),
  .ap_idle(PE_wrapper274_U0_ap_idle),
  .ap_ready(PE_wrapper274_U0_ap_ready),
  .fifo_cin_in_V_V_dout(fifo_cin_PE_10_4_V_V_dout),
  .fifo_cin_in_V_V_empty_n(fifo_cin_PE_10_4_V_V_empty_n),
  .fifo_cin_in_V_V_read(PE_wrapper274_U0_fifo_cin_in_V_V_read),
  .fifo_cin_out_V_V_din(PE_wrapper274_U0_fifo_cin_out_V_V_din),
  .fifo_cin_out_V_V_full_n(fifo_cin_PE_11_4_V_V_full_n),
  .fifo_cin_out_V_V_write(PE_wrapper274_U0_fifo_cin_out_V_V_write),
  .fifo_cout_drain_out_V_din(PE_wrapper274_U0_fifo_cout_drain_out_V_din),
  .fifo_cout_drain_out_V_full_n(fifo_cout_drain_PE_10_4_V_full_n),
  .fifo_cout_drain_out_V_write(PE_wrapper274_U0_fifo_cout_drain_out_V_write),
  .fifo_w_in_V_V_dout(fifo_w_PE_10_4_V_V_dout),
  .fifo_w_in_V_V_empty_n(fifo_w_PE_10_4_V_V_empty_n),
  .fifo_w_in_V_V_read(PE_wrapper274_U0_fifo_w_in_V_V_read),
  .fifo_w_out_V_V_din(PE_wrapper274_U0_fifo_w_out_V_V_din),
  .fifo_w_out_V_V_full_n(fifo_w_PE_10_5_V_V_full_n),
  .fifo_w_out_V_V_write(PE_wrapper274_U0_fifo_w_out_V_V_write)
);

(* keep_hierarchy = "yes" *)
kernel0_PE_wrapper286
PE_wrapper286_U0
(
  .ap_clk(ap_clk),
  .ap_rst(ap_rst_pipe),
  .ap_start(ap_start_pipe),
  .ap_done(PE_wrapper286_U0_ap_done),
  .ap_continue(1'b1),
  .ap_idle(PE_wrapper286_U0_ap_idle),
  .ap_ready(PE_wrapper286_U0_ap_ready),
  .fifo_cin_in_V_V_dout(fifo_cin_PE_11_4_V_V_dout),
  .fifo_cin_in_V_V_empty_n(fifo_cin_PE_11_4_V_V_empty_n),
  .fifo_cin_in_V_V_read(PE_wrapper286_U0_fifo_cin_in_V_V_read),
  .fifo_cin_out_V_V_din(PE_wrapper286_U0_fifo_cin_out_V_V_din),
  .fifo_cin_out_V_V_full_n(fifo_cin_PE_12_4_V_V_full_n),
  .fifo_cin_out_V_V_write(PE_wrapper286_U0_fifo_cin_out_V_V_write),
  .fifo_cout_drain_out_V_din(PE_wrapper286_U0_fifo_cout_drain_out_V_din),
  .fifo_cout_drain_out_V_full_n(fifo_cout_drain_PE_11_4_V_full_n),
  .fifo_cout_drain_out_V_write(PE_wrapper286_U0_fifo_cout_drain_out_V_write),
  .fifo_w_in_V_V_dout(fifo_w_PE_11_4_V_V_dout),
  .fifo_w_in_V_V_empty_n(fifo_w_PE_11_4_V_V_empty_n),
  .fifo_w_in_V_V_read(PE_wrapper286_U0_fifo_w_in_V_V_read),
  .fifo_w_out_V_V_din(PE_wrapper286_U0_fifo_w_out_V_V_din),
  .fifo_w_out_V_V_full_n(fifo_w_PE_11_5_V_V_full_n),
  .fifo_w_out_V_V_write(PE_wrapper286_U0_fifo_w_out_V_V_write)
);

(* keep_hierarchy = "yes" *)
kernel0_PE_wrapper318
PE_wrapper318_U0
(
  .ap_clk(ap_clk),
  .ap_rst(ap_rst_pipe),
  .ap_start(ap_start_pipe),
  .ap_done(PE_wrapper318_U0_ap_done),
  .ap_continue(1'b1),
  .ap_idle(PE_wrapper318_U0_ap_idle),
  .ap_ready(PE_wrapper318_U0_ap_ready),
  .fifo_cin_in_V_V_dout(fifo_cin_PE_14_0_V_V_dout),
  .fifo_cin_in_V_V_empty_n(fifo_cin_PE_14_0_V_V_empty_n),
  .fifo_cin_in_V_V_read(PE_wrapper318_U0_fifo_cin_in_V_V_read),
  .fifo_cin_out_V_V_din(PE_wrapper318_U0_fifo_cin_out_V_V_din),
  .fifo_cin_out_V_V_full_n(fifo_cin_PE_15_0_V_V_full_n),
  .fifo_cin_out_V_V_write(PE_wrapper318_U0_fifo_cin_out_V_V_write),
  .fifo_cout_drain_out_V_din(PE_wrapper318_U0_fifo_cout_drain_out_V_din),
  .fifo_cout_drain_out_V_full_n(fifo_cout_drain_PE_14_0_V_full_n),
  .fifo_cout_drain_out_V_write(PE_wrapper318_U0_fifo_cout_drain_out_V_write),
  .fifo_w_in_V_V_dout(fifo_w_PE_14_0_V_V_dout),
  .fifo_w_in_V_V_empty_n(fifo_w_PE_14_0_V_V_empty_n),
  .fifo_w_in_V_V_read(PE_wrapper318_U0_fifo_w_in_V_V_read),
  .fifo_w_out_V_V_din(PE_wrapper318_U0_fifo_w_out_V_V_din),
  .fifo_w_out_V_V_full_n(fifo_w_PE_14_1_V_V_full_n),
  .fifo_w_out_V_V_write(PE_wrapper318_U0_fifo_w_out_V_V_write)
);

(* keep_hierarchy = "yes" *)
kernel0_PE_wrapper320
PE_wrapper320_U0
(
  .ap_clk(ap_clk),
  .ap_rst(ap_rst_pipe),
  .ap_start(ap_start_pipe),
  .ap_done(PE_wrapper320_U0_ap_done),
  .ap_continue(1'b1),
  .ap_idle(PE_wrapper320_U0_ap_idle),
  .ap_ready(PE_wrapper320_U0_ap_ready),
  .fifo_cin_in_V_V_dout(fifo_cin_PE_14_2_V_V_dout),
  .fifo_cin_in_V_V_empty_n(fifo_cin_PE_14_2_V_V_empty_n),
  .fifo_cin_in_V_V_read(PE_wrapper320_U0_fifo_cin_in_V_V_read),
  .fifo_cin_out_V_V_din(PE_wrapper320_U0_fifo_cin_out_V_V_din),
  .fifo_cin_out_V_V_full_n(fifo_cin_PE_15_2_V_V_full_n),
  .fifo_cin_out_V_V_write(PE_wrapper320_U0_fifo_cin_out_V_V_write),
  .fifo_cout_drain_out_V_din(PE_wrapper320_U0_fifo_cout_drain_out_V_din),
  .fifo_cout_drain_out_V_full_n(fifo_cout_drain_PE_14_2_V_full_n),
  .fifo_cout_drain_out_V_write(PE_wrapper320_U0_fifo_cout_drain_out_V_write),
  .fifo_w_in_V_V_dout(fifo_w_PE_14_2_V_V_dout),
  .fifo_w_in_V_V_empty_n(fifo_w_PE_14_2_V_V_empty_n),
  .fifo_w_in_V_V_read(PE_wrapper320_U0_fifo_w_in_V_V_read),
  .fifo_w_out_V_V_din(PE_wrapper320_U0_fifo_w_out_V_V_din),
  .fifo_w_out_V_V_full_n(fifo_w_PE_14_3_V_V_full_n),
  .fifo_w_out_V_V_write(PE_wrapper320_U0_fifo_w_out_V_V_write)
);

(* keep_hierarchy = "yes" *)
kernel0_PE_wrapper321
PE_wrapper321_U0
(
  .ap_clk(ap_clk),
  .ap_rst(ap_rst_pipe),
  .ap_start(ap_start_pipe),
  .ap_done(PE_wrapper321_U0_ap_done),
  .ap_continue(1'b1),
  .ap_idle(PE_wrapper321_U0_ap_idle),
  .ap_ready(PE_wrapper321_U0_ap_ready),
  .fifo_cin_in_V_V_dout(fifo_cin_PE_14_3_V_V_dout),
  .fifo_cin_in_V_V_empty_n(fifo_cin_PE_14_3_V_V_empty_n),
  .fifo_cin_in_V_V_read(PE_wrapper321_U0_fifo_cin_in_V_V_read),
  .fifo_cin_out_V_V_din(PE_wrapper321_U0_fifo_cin_out_V_V_din),
  .fifo_cin_out_V_V_full_n(fifo_cin_PE_15_3_V_V_full_n),
  .fifo_cin_out_V_V_write(PE_wrapper321_U0_fifo_cin_out_V_V_write),
  .fifo_cout_drain_out_V_din(PE_wrapper321_U0_fifo_cout_drain_out_V_din),
  .fifo_cout_drain_out_V_full_n(fifo_cout_drain_PE_14_3_V_full_n),
  .fifo_cout_drain_out_V_write(PE_wrapper321_U0_fifo_cout_drain_out_V_write),
  .fifo_w_in_V_V_dout(fifo_w_PE_14_3_V_V_dout),
  .fifo_w_in_V_V_empty_n(fifo_w_PE_14_3_V_V_empty_n),
  .fifo_w_in_V_V_read(PE_wrapper321_U0_fifo_w_in_V_V_read),
  .fifo_w_out_V_V_din(PE_wrapper321_U0_fifo_w_out_V_V_din),
  .fifo_w_out_V_V_full_n(fifo_w_PE_14_4_V_V_full_n),
  .fifo_w_out_V_V_write(PE_wrapper321_U0_fifo_w_out_V_V_write)
);

(* keep_hierarchy = "yes" *)
kernel0_PE_wrapper330
PE_wrapper330_U0
(
  .ap_clk(ap_clk),
  .ap_rst(ap_rst_pipe),
  .ap_start(ap_start_pipe),
  .ap_done(PE_wrapper330_U0_ap_done),
  .ap_continue(1'b1),
  .ap_idle(PE_wrapper330_U0_ap_idle),
  .ap_ready(PE_wrapper330_U0_ap_ready),
  .fifo_cin_in_V_V_dout(fifo_cin_PE_15_0_V_V_dout),
  .fifo_cin_in_V_V_empty_n(fifo_cin_PE_15_0_V_V_empty_n),
  .fifo_cin_in_V_V_read(PE_wrapper330_U0_fifo_cin_in_V_V_read),
  .fifo_cin_out_V_V_din(PE_wrapper330_U0_fifo_cin_out_V_V_din),
  .fifo_cin_out_V_V_full_n(fifo_cin_PE_16_0_V_V_full_n),
  .fifo_cin_out_V_V_write(PE_wrapper330_U0_fifo_cin_out_V_V_write),
  .fifo_cout_drain_out_V_din(PE_wrapper330_U0_fifo_cout_drain_out_V_din),
  .fifo_cout_drain_out_V_full_n(fifo_cout_drain_PE_15_0_V_full_n),
  .fifo_cout_drain_out_V_write(PE_wrapper330_U0_fifo_cout_drain_out_V_write),
  .fifo_w_in_V_V_dout(fifo_w_PE_15_0_V_V_dout),
  .fifo_w_in_V_V_empty_n(fifo_w_PE_15_0_V_V_empty_n),
  .fifo_w_in_V_V_read(PE_wrapper330_U0_fifo_w_in_V_V_read),
  .fifo_w_out_V_V_din(PE_wrapper330_U0_fifo_w_out_V_V_din),
  .fifo_w_out_V_V_full_n(fifo_w_PE_15_1_V_V_full_n),
  .fifo_w_out_V_V_write(PE_wrapper330_U0_fifo_w_out_V_V_write)
);

(* keep_hierarchy = "yes" *)
kernel0_cout_drain_IO_L1_out_wrapper384
cout_drain_IO_L1_out_wrapper384_U0
(
  .ap_clk(ap_clk),
  .ap_rst(ap_rst_pipe),
  .ap_start(ap_start_pipe),
  .ap_done(cout_drain_IO_L1_out_wrapper384_U0_ap_done),
  .ap_continue(1'b1),
  .ap_idle(cout_drain_IO_L1_out_wrapper384_U0_ap_idle),
  .ap_ready(cout_drain_IO_L1_out_wrapper384_U0_ap_ready),
  .fifo_cout_drain_in_V_V_dout(fifo_cout_drain_cout_drain_IO_L1_out_1_15_V_V_dout),
  .fifo_cout_drain_in_V_V_empty_n(fifo_cout_drain_cout_drain_IO_L1_out_1_15_V_V_empty_n),
  .fifo_cout_drain_in_V_V_read(cout_drain_IO_L1_out_wrapper384_U0_fifo_cout_drain_in_V_V_read),
  .fifo_cout_drain_out_V_V_din(cout_drain_IO_L1_out_wrapper384_U0_fifo_cout_drain_out_V_V_din),
  .fifo_cout_drain_out_V_V_full_n(fifo_cout_drain_cout_drain_IO_L1_out_1_14_V_V_full_n),
  .fifo_cout_drain_out_V_V_write(cout_drain_IO_L1_out_wrapper384_U0_fifo_cout_drain_out_V_V_write),
  .fifo_cout_drain_local_in_V_dout(fifo_cout_drain_PE_14_1_V_dout),
  .fifo_cout_drain_local_in_V_empty_n(fifo_cout_drain_PE_14_1_V_empty_n),
  .fifo_cout_drain_local_in_V_read(cout_drain_IO_L1_out_wrapper384_U0_fifo_cout_drain_local_in_V_read)
);

(* keep_hierarchy = "yes" *)
kernel0_cout_drain_IO_L1_out_wrapper402
cout_drain_IO_L1_out_wrapper402_U0
(
  .ap_clk(ap_clk),
  .ap_rst(ap_rst_pipe),
  .ap_start(ap_start_pipe),
  .ap_done(cout_drain_IO_L1_out_wrapper402_U0_ap_done),
  .ap_continue(1'b1),
  .ap_idle(cout_drain_IO_L1_out_wrapper402_U0_ap_idle),
  .ap_ready(cout_drain_IO_L1_out_wrapper402_U0_ap_ready),
  .fifo_cout_drain_in_V_V_dout(fifo_cout_drain_cout_drain_IO_L1_out_2_13_V_V_dout),
  .fifo_cout_drain_in_V_V_empty_n(fifo_cout_drain_cout_drain_IO_L1_out_2_13_V_V_empty_n),
  .fifo_cout_drain_in_V_V_read(cout_drain_IO_L1_out_wrapper402_U0_fifo_cout_drain_in_V_V_read),
  .fifo_cout_drain_out_V_V_din(cout_drain_IO_L1_out_wrapper402_U0_fifo_cout_drain_out_V_V_din),
  .fifo_cout_drain_out_V_V_full_n(fifo_cout_drain_cout_drain_IO_L1_out_2_12_V_V_full_n),
  .fifo_cout_drain_out_V_V_write(cout_drain_IO_L1_out_wrapper402_U0_fifo_cout_drain_out_V_V_write),
  .fifo_cout_drain_local_in_V_dout(fifo_cout_drain_PE_12_2_V_dout),
  .fifo_cout_drain_local_in_V_empty_n(fifo_cout_drain_PE_12_2_V_empty_n),
  .fifo_cout_drain_local_in_V_read(cout_drain_IO_L1_out_wrapper402_U0_fifo_cout_drain_local_in_V_read)
);

(* keep_hierarchy = "yes" *)
kernel0_cout_drain_IO_L1_out_wrapper416
cout_drain_IO_L1_out_wrapper416_U0
(
  .ap_clk(ap_clk),
  .ap_rst(ap_rst_pipe),
  .ap_start(ap_start_pipe),
  .ap_done(cout_drain_IO_L1_out_wrapper416_U0_ap_done),
  .ap_continue(1'b1),
  .ap_idle(cout_drain_IO_L1_out_wrapper416_U0_ap_idle),
  .ap_ready(cout_drain_IO_L1_out_wrapper416_U0_ap_ready),
  .fifo_cout_drain_in_V_V_dout(fifo_cout_drain_cout_drain_IO_L1_out_3_15_V_V_dout),
  .fifo_cout_drain_in_V_V_empty_n(fifo_cout_drain_cout_drain_IO_L1_out_3_15_V_V_empty_n),
  .fifo_cout_drain_in_V_V_read(cout_drain_IO_L1_out_wrapper416_U0_fifo_cout_drain_in_V_V_read),
  .fifo_cout_drain_out_V_V_din(cout_drain_IO_L1_out_wrapper416_U0_fifo_cout_drain_out_V_V_din),
  .fifo_cout_drain_out_V_V_full_n(fifo_cout_drain_cout_drain_IO_L1_out_3_14_V_V_full_n),
  .fifo_cout_drain_out_V_V_write(cout_drain_IO_L1_out_wrapper416_U0_fifo_cout_drain_out_V_V_write),
  .fifo_cout_drain_local_in_V_dout(fifo_cout_drain_PE_14_3_V_dout),
  .fifo_cout_drain_local_in_V_empty_n(fifo_cout_drain_PE_14_3_V_empty_n),
  .fifo_cout_drain_local_in_V_read(cout_drain_IO_L1_out_wrapper416_U0_fifo_cout_drain_local_in_V_read)
);

(* keep_hierarchy = "yes" *)
kernel0_cout_drain_IO_L1_out_wrapper419
cout_drain_IO_L1_out_wrapper419_U0
(
  .ap_clk(ap_clk),
  .ap_rst(ap_rst_pipe),
  .ap_start(ap_start_pipe),
  .ap_done(cout_drain_IO_L1_out_wrapper419_U0_ap_done),
  .ap_continue(1'b1),
  .ap_idle(cout_drain_IO_L1_out_wrapper419_U0_ap_idle),
  .ap_ready(cout_drain_IO_L1_out_wrapper419_U0_ap_ready),
  .fifo_cout_drain_in_V_V_dout(fifo_cout_drain_cout_drain_IO_L1_out_3_12_V_V_dout),
  .fifo_cout_drain_in_V_V_empty_n(fifo_cout_drain_cout_drain_IO_L1_out_3_12_V_V_empty_n),
  .fifo_cout_drain_in_V_V_read(cout_drain_IO_L1_out_wrapper419_U0_fifo_cout_drain_in_V_V_read),
  .fifo_cout_drain_out_V_V_din(cout_drain_IO_L1_out_wrapper419_U0_fifo_cout_drain_out_V_V_din),
  .fifo_cout_drain_out_V_V_full_n(fifo_cout_drain_cout_drain_IO_L1_out_3_11_V_V_full_n),
  .fifo_cout_drain_out_V_V_write(cout_drain_IO_L1_out_wrapper419_U0_fifo_cout_drain_out_V_V_write),
  .fifo_cout_drain_local_in_V_dout(fifo_cout_drain_PE_11_3_V_dout),
  .fifo_cout_drain_local_in_V_empty_n(fifo_cout_drain_PE_11_3_V_empty_n),
  .fifo_cout_drain_local_in_V_read(cout_drain_IO_L1_out_wrapper419_U0_fifo_cout_drain_local_in_V_read)
);

(* keep_hierarchy = "yes" *)
kernel0_cout_drain_IO_L1_out_boundary_wrapper431
cout_drain_IO_L1_out_boundary_wrapper431_U0
(
  .ap_clk(ap_clk),
  .ap_rst(ap_rst_pipe),
  .ap_start(ap_start_pipe),
  .ap_done(cout_drain_IO_L1_out_boundary_wrapper431_U0_ap_done),
  .ap_continue(1'b1),
  .ap_idle(cout_drain_IO_L1_out_boundary_wrapper431_U0_ap_idle),
  .ap_ready(cout_drain_IO_L1_out_boundary_wrapper431_U0_ap_ready),
  .fifo_cout_drain_out_V_V_din(cout_drain_IO_L1_out_boundary_wrapper431_U0_fifo_cout_drain_out_V_V_din),
  .fifo_cout_drain_out_V_V_full_n(fifo_cout_drain_cout_drain_IO_L1_out_4_15_V_V_full_n),
  .fifo_cout_drain_out_V_V_write(cout_drain_IO_L1_out_boundary_wrapper431_U0_fifo_cout_drain_out_V_V_write),
  .fifo_cout_drain_local_in_V_dout(fifo_cout_drain_PE_15_4_V_dout),
  .fifo_cout_drain_local_in_V_empty_n(fifo_cout_drain_PE_15_4_V_empty_n),
  .fifo_cout_drain_local_in_V_read(cout_drain_IO_L1_out_boundary_wrapper431_U0_fifo_cout_drain_local_in_V_read)
);

(* keep_hierarchy = "yes" *)
kernel0_cout_drain_IO_L1_out_wrapper432
cout_drain_IO_L1_out_wrapper432_U0
(
  .ap_clk(ap_clk),
  .ap_rst(ap_rst_pipe),
  .ap_start(ap_start_pipe),
  .ap_done(cout_drain_IO_L1_out_wrapper432_U0_ap_done),
  .ap_continue(1'b1),
  .ap_idle(cout_drain_IO_L1_out_wrapper432_U0_ap_idle),
  .ap_ready(cout_drain_IO_L1_out_wrapper432_U0_ap_ready),
  .fifo_cout_drain_in_V_V_dout(fifo_cout_drain_cout_drain_IO_L1_out_4_15_V_V_dout),
  .fifo_cout_drain_in_V_V_empty_n(fifo_cout_drain_cout_drain_IO_L1_out_4_15_V_V_empty_n),
  .fifo_cout_drain_in_V_V_read(cout_drain_IO_L1_out_wrapper432_U0_fifo_cout_drain_in_V_V_read),
  .fifo_cout_drain_out_V_V_din(cout_drain_IO_L1_out_wrapper432_U0_fifo_cout_drain_out_V_V_din),
  .fifo_cout_drain_out_V_V_full_n(fifo_cout_drain_cout_drain_IO_L1_out_4_14_V_V_full_n),
  .fifo_cout_drain_out_V_V_write(cout_drain_IO_L1_out_wrapper432_U0_fifo_cout_drain_out_V_V_write),
  .fifo_cout_drain_local_in_V_dout(fifo_cout_drain_PE_14_4_V_dout),
  .fifo_cout_drain_local_in_V_empty_n(fifo_cout_drain_PE_14_4_V_empty_n),
  .fifo_cout_drain_local_in_V_read(cout_drain_IO_L1_out_wrapper432_U0_fifo_cout_drain_local_in_V_read)
);

(* keep_hierarchy = "yes" *)
kernel0_cout_drain_IO_L1_out_wrapper434
cout_drain_IO_L1_out_wrapper434_U0
(
  .ap_clk(ap_clk),
  .ap_rst(ap_rst_pipe),
  .ap_start(ap_start_pipe),
  .ap_done(cout_drain_IO_L1_out_wrapper434_U0_ap_done),
  .ap_continue(1'b1),
  .ap_idle(cout_drain_IO_L1_out_wrapper434_U0_ap_idle),
  .ap_ready(cout_drain_IO_L1_out_wrapper434_U0_ap_ready),
  .fifo_cout_drain_in_V_V_dout(fifo_cout_drain_cout_drain_IO_L1_out_4_13_V_V_dout),
  .fifo_cout_drain_in_V_V_empty_n(fifo_cout_drain_cout_drain_IO_L1_out_4_13_V_V_empty_n),
  .fifo_cout_drain_in_V_V_read(cout_drain_IO_L1_out_wrapper434_U0_fifo_cout_drain_in_V_V_read),
  .fifo_cout_drain_out_V_V_din(cout_drain_IO_L1_out_wrapper434_U0_fifo_cout_drain_out_V_V_din),
  .fifo_cout_drain_out_V_V_full_n(fifo_cout_drain_cout_drain_IO_L1_out_4_12_V_V_full_n),
  .fifo_cout_drain_out_V_V_write(cout_drain_IO_L1_out_wrapper434_U0_fifo_cout_drain_out_V_V_write),
  .fifo_cout_drain_local_in_V_dout(fifo_cout_drain_PE_12_4_V_dout),
  .fifo_cout_drain_local_in_V_empty_n(fifo_cout_drain_PE_12_4_V_empty_n),
  .fifo_cout_drain_local_in_V_read(cout_drain_IO_L1_out_wrapper434_U0_fifo_cout_drain_local_in_V_read)
);

(* keep_hierarchy = "yes" *)
fifo_almost_full
#(
  .DATA_WIDTH(256),
  .DEPTH(3),
  .ADDR_WIDTH(9),
  .GRACE_PERIOD(1)
)
fifo_cin_PE_11_4_V_V_U
(
  .clk(ap_clk),
  .reset(ap_rst_n_inv),
  .if_read_ce(1'b1),
  .if_write_ce(1'b1),
  .if_din(PE_wrapper274_U0_fifo_cin_out_V_V_din),
  .if_full_n(fifo_cin_PE_11_4_V_V_full_n),
  .if_write(PE_wrapper274_U0_fifo_cin_out_V_V_write),
  .if_dout(fifo_cin_PE_11_4_V_V_dout),
  .if_empty_n(fifo_cin_PE_11_4_V_V_empty_n),
  .if_read(PE_wrapper286_U0_fifo_cin_in_V_V_read)
);

(* keep_hierarchy = "yes" *)
fifo_almost_full
#(
  .DATA_WIDTH(32),
  .DEPTH(9),
  .ADDR_WIDTH(6),
  .GRACE_PERIOD(1)
)
fifo_cout_drain_PE_14_3_V_U
(
  .clk(ap_clk),
  .reset(ap_rst_n_inv),
  .if_read_ce(1'b1),
  .if_write_ce(1'b1),
  .if_din(PE_wrapper321_U0_fifo_cout_drain_out_V_din),
  .if_full_n(fifo_cout_drain_PE_14_3_V_full_n),
  .if_write(PE_wrapper321_U0_fifo_cout_drain_out_V_write),
  .if_dout(fifo_cout_drain_PE_14_3_V_dout),
  .if_empty_n(fifo_cout_drain_PE_14_3_V_empty_n),
  .if_read(cout_drain_IO_L1_out_wrapper416_U0_fifo_cout_drain_local_in_V_read)
);

(* keep_hierarchy = "yes" *)
fifo_almost_full
#(
  .DATA_WIDTH(256),
  .DEPTH(5),
  .ADDR_WIDTH(9),
  .GRACE_PERIOD(1)
)
fifo_w_PE_14_3_V_V_U
(
  .clk(ap_clk),
  .reset(ap_rst_n_inv),
  .if_read_ce(1'b1),
  .if_write_ce(1'b1),
  .if_din(PE_wrapper320_U0_fifo_w_out_V_V_din),
  .if_full_n(fifo_w_PE_14_3_V_V_full_n),
  .if_write(PE_wrapper320_U0_fifo_w_out_V_V_write),
  .if_dout(fifo_w_PE_14_3_V_V_dout),
  .if_empty_n(fifo_w_PE_14_3_V_V_empty_n),
  .if_read(PE_wrapper321_U0_fifo_w_in_V_V_read)
);

(* keep_hierarchy = "yes" *)
fifo_almost_full
#(
  .DATA_WIDTH(256),
  .DEPTH(3),
  .ADDR_WIDTH(9),
  .GRACE_PERIOD(1)
)
fifo_cin_PE_15_0_V_V_U
(
  .clk(ap_clk),
  .reset(ap_rst_n_inv),
  .if_read_ce(1'b1),
  .if_write_ce(1'b1),
  .if_din(PE_wrapper318_U0_fifo_cin_out_V_V_din),
  .if_full_n(fifo_cin_PE_15_0_V_V_full_n),
  .if_write(PE_wrapper318_U0_fifo_cin_out_V_V_write),
  .if_dout(fifo_cin_PE_15_0_V_V_dout),
  .if_empty_n(fifo_cin_PE_15_0_V_V_empty_n),
  .if_read(PE_wrapper330_U0_fifo_cin_in_V_V_read)
);

(* keep_hierarchy = "yes" *)
fifo_almost_full
#(
  .DATA_WIDTH(64),
  .DEPTH(3),
  .ADDR_WIDTH(7),
  .GRACE_PERIOD(1)
)
fifo_cout_drain_cout_drain_IO_L1_out_4_15_V_V_U
(
  .clk(ap_clk),
  .reset(ap_rst_n_inv),
  .if_read_ce(1'b1),
  .if_write_ce(1'b1),
  .if_din(cout_drain_IO_L1_out_boundary_wrapper431_U0_fifo_cout_drain_out_V_V_din),
  .if_full_n(fifo_cout_drain_cout_drain_IO_L1_out_4_15_V_V_full_n),
  .if_write(cout_drain_IO_L1_out_boundary_wrapper431_U0_fifo_cout_drain_out_V_V_write),
  .if_dout(fifo_cout_drain_cout_drain_IO_L1_out_4_15_V_V_dout),
  .if_empty_n(fifo_cout_drain_cout_drain_IO_L1_out_4_15_V_V_empty_n),
  .if_read(cout_drain_IO_L1_out_wrapper432_U0_fifo_cout_drain_in_V_V_read)
);

(* keep_hierarchy = "yes" *)
fifo_almost_full
#(
  .DATA_WIDTH(256),
  .DEPTH(5),
  .ADDR_WIDTH(9),
  .GRACE_PERIOD(1)
)
fifo_w_PE_14_0_V_V_U
(
  .clk(ap_clk),
  .reset(ap_rst_n_inv),
  .if_read_ce(1'b1),
  .if_write_ce(1'b1),
  .if_din(w_IO_L2_in149_U0_fifo_w_local_out_V_V_din),
  .if_full_n(fifo_w_PE_14_0_V_V_full_n),
  .if_write(w_IO_L2_in149_U0_fifo_w_local_out_V_V_write),
  .if_dout(fifo_w_PE_14_0_V_V_dout),
  .if_empty_n(fifo_w_PE_14_0_V_V_empty_n),
  .if_read(PE_wrapper318_U0_fifo_w_in_V_V_read)
);

(* keep_hierarchy = "yes" *)
fifo_almost_full
#(
  .DATA_WIDTH(64),
  .DEPTH(4),
  .ADDR_WIDTH(7),
  .GRACE_PERIOD(3)
)
fifo_cout_drain_cout_drain_IO_L1_out_4_13_V_V_U
(
  .clk(ap_clk),
  .reset(ap_rst_n_inv),
  .if_read_ce(1'b1),
  .if_write_ce(1'b1),
  .if_din(cout_drain_IO_L1_out_wrapper433_U0_fifo_cout_drain_out_V_V_din),
  .if_full_n(fifo_cout_drain_cout_drain_IO_L1_out_4_13_V_V_full_n),
  .if_write(cout_drain_IO_L1_out_wrapper433_U0_fifo_cout_drain_out_V_V_write),
  .if_dout(fifo_cout_drain_cout_drain_IO_L1_out_4_13_V_V_dout),
  .if_empty_n(fifo_cout_drain_cout_drain_IO_L1_out_4_13_V_V_empty_n),
  .if_read(cout_drain_IO_L1_out_wrapper434_U0_fifo_cout_drain_in_V_V_read)
);

(* keep_hierarchy = "yes" *)
fifo_almost_full
#(
  .DATA_WIDTH(256),
  .DEPTH(5),
  .ADDR_WIDTH(9),
  .GRACE_PERIOD(5)
)
fifo_cin_PE_14_3_V_V_U
(
  .clk(ap_clk),
  .reset(ap_rst_n_inv),
  .if_read_ce(1'b1),
  .if_write_ce(1'b1),
  .if_din(PE_wrapper309_U0_fifo_cin_out_V_V_din),
  .if_full_n(fifo_cin_PE_14_3_V_V_full_n),
  .if_write(PE_wrapper309_U0_fifo_cin_out_V_V_write),
  .if_dout(fifo_cin_PE_14_3_V_V_dout),
  .if_empty_n(fifo_cin_PE_14_3_V_V_empty_n),
  .if_read(PE_wrapper321_U0_fifo_cin_in_V_V_read)
);

(* keep_hierarchy = "yes" *)
fifo_almost_full
#(
  .DATA_WIDTH(256),
  .DEPTH(5),
  .ADDR_WIDTH(9),
  .GRACE_PERIOD(5)
)
fifo_cin_PE_6_4_V_V_U
(
  .clk(ap_clk),
  .reset(ap_rst_n_inv),
  .if_read_ce(1'b1),
  .if_write_ce(1'b1),
  .if_din(PE_wrapper214_U0_fifo_cin_out_V_V_din),
  .if_full_n(fifo_cin_PE_6_4_V_V_full_n),
  .if_write(PE_wrapper214_U0_fifo_cin_out_V_V_write),
  .if_dout(fifo_cin_PE_6_4_V_V_dout),
  .if_empty_n(fifo_cin_PE_6_4_V_V_empty_n),
  .if_read(PE_wrapper226_U0_fifo_cin_in_V_V_read)
);

(* keep_hierarchy = "yes" *)
fifo_almost_full
#(
  .DATA_WIDTH(256),
  .DEPTH(4),
  .ADDR_WIDTH(9),
  .GRACE_PERIOD(3)
)
fifo_w_w_IO_L2_in_14_V_V_U
(
  .clk(ap_clk),
  .reset(ap_rst_n_inv),
  .if_read_ce(1'b1),
  .if_write_ce(1'b1),
  .if_din(w_IO_L2_in148_U0_fifo_w_out_V_V_din),
  .if_full_n(fifo_w_w_IO_L2_in_14_V_V_full_n),
  .if_write(w_IO_L2_in148_U0_fifo_w_out_V_V_write),
  .if_dout(fifo_w_w_IO_L2_in_14_V_V_dout),
  .if_empty_n(fifo_w_w_IO_L2_in_14_V_V_empty_n),
  .if_read(w_IO_L2_in149_U0_fifo_w_in_V_V_read)
);

(* keep_hierarchy = "yes" *)
fifo_almost_full
#(
  .DATA_WIDTH(64),
  .DEPTH(5),
  .ADDR_WIDTH(7),
  .GRACE_PERIOD(5)
)
fifo_cout_drain_cout_drain_IO_L1_out_3_12_V_V_U
(
  .clk(ap_clk),
  .reset(ap_rst_n_inv),
  .if_read_ce(1'b1),
  .if_write_ce(1'b1),
  .if_din(cout_drain_IO_L1_out_wrapper418_U0_fifo_cout_drain_out_V_V_din),
  .if_full_n(fifo_cout_drain_cout_drain_IO_L1_out_3_12_V_V_full_n),
  .if_write(cout_drain_IO_L1_out_wrapper418_U0_fifo_cout_drain_out_V_V_write),
  .if_dout(fifo_cout_drain_cout_drain_IO_L1_out_3_12_V_V_dout),
  .if_empty_n(fifo_cout_drain_cout_drain_IO_L1_out_3_12_V_V_empty_n),
  .if_read(cout_drain_IO_L1_out_wrapper419_U0_fifo_cout_drain_in_V_V_read)
);

(* keep_hierarchy = "yes" *)
fifo_almost_full
#(
  .DATA_WIDTH(256),
  .DEPTH(5),
  .ADDR_WIDTH(9),
  .GRACE_PERIOD(5)
)
fifo_w_PE_6_4_V_V_U
(
  .clk(ap_clk),
  .reset(ap_rst_n_inv),
  .if_read_ce(1'b1),
  .if_write_ce(1'b1),
  .if_din(PE_wrapper225_U0_fifo_w_out_V_V_din),
  .if_full_n(fifo_w_PE_6_4_V_V_full_n),
  .if_write(PE_wrapper225_U0_fifo_w_out_V_V_write),
  .if_dout(fifo_w_PE_6_4_V_V_dout),
  .if_empty_n(fifo_w_PE_6_4_V_V_empty_n),
  .if_read(PE_wrapper226_U0_fifo_w_in_V_V_read)
);

(* keep_hierarchy = "yes" *)
fifo_almost_full
#(
  .DATA_WIDTH(256),
  .DEPTH(5),
  .ADDR_WIDTH(9),
  .GRACE_PERIOD(5)
)
fifo_w_PE_11_4_V_V_U
(
  .clk(ap_clk),
  .reset(ap_rst_n_inv),
  .if_read_ce(1'b1),
  .if_write_ce(1'b1),
  .if_din(PE_wrapper285_U0_fifo_w_out_V_V_din),
  .if_full_n(fifo_w_PE_11_4_V_V_full_n),
  .if_write(PE_wrapper285_U0_fifo_w_out_V_V_write),
  .if_dout(fifo_w_PE_11_4_V_V_dout),
  .if_empty_n(fifo_w_PE_11_4_V_V_empty_n),
  .if_read(PE_wrapper286_U0_fifo_w_in_V_V_read)
);

(* keep_hierarchy = "yes" *)
fifo_almost_full
#(
  .DATA_WIDTH(256),
  .DEPTH(4),
  .ADDR_WIDTH(9),
  .GRACE_PERIOD(3)
)
fifo_w_PE_15_0_V_V_U
(
  .clk(ap_clk),
  .reset(ap_rst_n_inv),
  .if_read_ce(1'b1),
  .if_write_ce(1'b1),
  .if_din(w_IO_L2_in_boundary_U0_fifo_w_local_out_V_V_din),
  .if_full_n(fifo_w_PE_15_0_V_V_full_n),
  .if_write(w_IO_L2_in_boundary_U0_fifo_w_local_out_V_V_write),
  .if_dout(fifo_w_PE_15_0_V_V_dout),
  .if_empty_n(fifo_w_PE_15_0_V_V_empty_n),
  .if_read(PE_wrapper330_U0_fifo_w_in_V_V_read)
);

(* keep_hierarchy = "yes" *)
fifo_almost_full
#(
  .DATA_WIDTH(256),
  .DEPTH(6),
  .ADDR_WIDTH(9),
  .GRACE_PERIOD(3)
)
fifo_w_PE_10_4_V_V_U
(
  .clk(ap_clk),
  .reset(ap_rst_n_inv),
  .if_read_ce(1'b1),
  .if_write_ce(1'b1),
  .if_din(PE_wrapper273_U0_fifo_w_out_V_V_din),
  .if_full_n(fifo_w_PE_10_4_V_V_full_n),
  .if_write(PE_wrapper273_U0_fifo_w_out_V_V_write),
  .if_dout(fifo_w_PE_10_4_V_V_dout),
  .if_empty_n(fifo_w_PE_10_4_V_V_empty_n),
  .if_read(PE_wrapper274_U0_fifo_w_in_V_V_read)
);

(* keep_hierarchy = "yes" *)
fifo_almost_full
#(
  .DATA_WIDTH(64),
  .DEPTH(4),
  .ADDR_WIDTH(7),
  .GRACE_PERIOD(3)
)
fifo_cout_drain_cout_drain_IO_L1_out_1_15_V_V_U
(
  .clk(ap_clk),
  .reset(ap_rst_n_inv),
  .if_read_ce(1'b1),
  .if_write_ce(1'b1),
  .if_din(cout_drain_IO_L1_out_boundary_wrapper383_U0_fifo_cout_drain_out_V_V_din),
  .if_full_n(fifo_cout_drain_cout_drain_IO_L1_out_1_15_V_V_full_n),
  .if_write(cout_drain_IO_L1_out_boundary_wrapper383_U0_fifo_cout_drain_out_V_V_write),
  .if_dout(fifo_cout_drain_cout_drain_IO_L1_out_1_15_V_V_dout),
  .if_empty_n(fifo_cout_drain_cout_drain_IO_L1_out_1_15_V_V_empty_n),
  .if_read(cout_drain_IO_L1_out_wrapper384_U0_fifo_cout_drain_in_V_V_read)
);

(* keep_hierarchy = "yes" *)
fifo_almost_full
#(
  .DATA_WIDTH(256),
  .DEPTH(5),
  .ADDR_WIDTH(9),
  .GRACE_PERIOD(5)
)
fifo_cin_PE_14_0_V_V_U
(
  .clk(ap_clk),
  .reset(ap_rst_n_inv),
  .if_read_ce(1'b1),
  .if_write_ce(1'b1),
  .if_din(PE_wrapper306_U0_fifo_cin_out_V_V_din),
  .if_full_n(fifo_cin_PE_14_0_V_V_full_n),
  .if_write(PE_wrapper306_U0_fifo_cin_out_V_V_write),
  .if_dout(fifo_cin_PE_14_0_V_V_dout),
  .if_empty_n(fifo_cin_PE_14_0_V_V_empty_n),
  .if_read(PE_wrapper318_U0_fifo_cin_in_V_V_read)
);

(* keep_hierarchy = "yes" *)
fifo_almost_full
#(
  .DATA_WIDTH(32),
  .DEPTH(23),
  .ADDR_WIDTH(6),
  .GRACE_PERIOD(5)
)
fifo_cout_drain_PE_11_3_V_U
(
  .clk(ap_clk),
  .reset(ap_rst_n_inv),
  .if_read_ce(1'b1),
  .if_write_ce(1'b1),
  .if_din(PE_wrapper285_U0_fifo_cout_drain_out_V_din),
  .if_full_n(fifo_cout_drain_PE_11_3_V_full_n),
  .if_write(PE_wrapper285_U0_fifo_cout_drain_out_V_write),
  .if_dout(fifo_cout_drain_PE_11_3_V_dout),
  .if_empty_n(fifo_cout_drain_PE_11_3_V_empty_n),
  .if_read(cout_drain_IO_L1_out_wrapper419_U0_fifo_cout_drain_local_in_V_read)
);

(* keep_hierarchy = "yes" *)
fifo_almost_full
#(
  .DATA_WIDTH(256),
  .DEPTH(4),
  .ADDR_WIDTH(9),
  .GRACE_PERIOD(3)
)
fifo_w_PE_14_2_V_V_U
(
  .clk(ap_clk),
  .reset(ap_rst_n_inv),
  .if_read_ce(1'b1),
  .if_write_ce(1'b1),
  .if_din(PE_wrapper319_U0_fifo_w_out_V_V_din),
  .if_full_n(fifo_w_PE_14_2_V_V_full_n),
  .if_write(PE_wrapper319_U0_fifo_w_out_V_V_write),
  .if_dout(fifo_w_PE_14_2_V_V_dout),
  .if_empty_n(fifo_w_PE_14_2_V_V_empty_n),
  .if_read(PE_wrapper320_U0_fifo_w_in_V_V_read)
);

(* keep_hierarchy = "yes" *)
fifo_almost_full
#(
  .DATA_WIDTH(256),
  .DEPTH(4),
  .ADDR_WIDTH(9),
  .GRACE_PERIOD(3)
)
fifo_cin_PE_14_2_V_V_U
(
  .clk(ap_clk),
  .reset(ap_rst_n_inv),
  .if_read_ce(1'b1),
  .if_write_ce(1'b1),
  .if_din(PE_wrapper308_U0_fifo_cin_out_V_V_din),
  .if_full_n(fifo_cin_PE_14_2_V_V_full_n),
  .if_write(PE_wrapper308_U0_fifo_cin_out_V_V_write),
  .if_dout(fifo_cin_PE_14_2_V_V_dout),
  .if_empty_n(fifo_cin_PE_14_2_V_V_empty_n),
  .if_read(PE_wrapper320_U0_fifo_cin_in_V_V_read)
);

(* keep_hierarchy = "yes" *)
fifo_almost_full
#(
  .DATA_WIDTH(32),
  .DEPTH(6),
  .ADDR_WIDTH(6),
  .GRACE_PERIOD(3)
)
fifo_cout_drain_PE_14_1_V_U
(
  .clk(ap_clk),
  .reset(ap_rst_n_inv),
  .if_read_ce(1'b1),
  .if_write_ce(1'b1),
  .if_din(PE_wrapper319_U0_fifo_cout_drain_out_V_din),
  .if_full_n(fifo_cout_drain_PE_14_1_V_full_n),
  .if_write(PE_wrapper319_U0_fifo_cout_drain_out_V_write),
  .if_dout(fifo_cout_drain_PE_14_1_V_dout),
  .if_empty_n(fifo_cout_drain_PE_14_1_V_empty_n),
  .if_read(cout_drain_IO_L1_out_wrapper384_U0_fifo_cout_drain_local_in_V_read)
);

(* keep_hierarchy = "yes" *)
fifo_almost_full
#(
  .DATA_WIDTH(32),
  .DEPTH(4),
  .ADDR_WIDTH(6),
  .GRACE_PERIOD(3)
)
fifo_cout_drain_PE_15_4_V_U
(
  .clk(ap_clk),
  .reset(ap_rst_n_inv),
  .if_read_ce(1'b1),
  .if_write_ce(1'b1),
  .if_din(PE_wrapper334_U0_fifo_cout_drain_out_V_din),
  .if_full_n(fifo_cout_drain_PE_15_4_V_full_n),
  .if_write(PE_wrapper334_U0_fifo_cout_drain_out_V_write),
  .if_dout(fifo_cout_drain_PE_15_4_V_dout),
  .if_empty_n(fifo_cout_drain_PE_15_4_V_empty_n),
  .if_read(cout_drain_IO_L1_out_boundary_wrapper431_U0_fifo_cout_drain_local_in_V_read)
);

(* keep_hierarchy = "yes" *)
fifo_almost_full
#(
  .DATA_WIDTH(64),
  .DEPTH(4),
  .ADDR_WIDTH(7),
  .GRACE_PERIOD(3)
)
fifo_cout_drain_cout_drain_IO_L1_out_3_15_V_V_U
(
  .clk(ap_clk),
  .reset(ap_rst_n_inv),
  .if_read_ce(1'b1),
  .if_write_ce(1'b1),
  .if_din(cout_drain_IO_L1_out_boundary_wrapper415_U0_fifo_cout_drain_out_V_V_din),
  .if_full_n(fifo_cout_drain_cout_drain_IO_L1_out_3_15_V_V_full_n),
  .if_write(cout_drain_IO_L1_out_boundary_wrapper415_U0_fifo_cout_drain_out_V_V_write),
  .if_dout(fifo_cout_drain_cout_drain_IO_L1_out_3_15_V_V_dout),
  .if_empty_n(fifo_cout_drain_cout_drain_IO_L1_out_3_15_V_V_empty_n),
  .if_read(cout_drain_IO_L1_out_wrapper416_U0_fifo_cout_drain_in_V_V_read)
);

(* keep_hierarchy = "yes" *)
fifo_almost_full
#(
  .DATA_WIDTH(256),
  .DEPTH(5),
  .ADDR_WIDTH(9),
  .GRACE_PERIOD(5)
)
fifo_cin_PE_10_4_V_V_U
(
  .clk(ap_clk),
  .reset(ap_rst_n_inv),
  .if_read_ce(1'b1),
  .if_write_ce(1'b1),
  .if_din(PE_wrapper262_U0_fifo_cin_out_V_V_din),
  .if_full_n(fifo_cin_PE_10_4_V_V_full_n),
  .if_write(PE_wrapper262_U0_fifo_cin_out_V_V_write),
  .if_dout(fifo_cin_PE_10_4_V_V_dout),
  .if_empty_n(fifo_cin_PE_10_4_V_V_empty_n),
  .if_read(PE_wrapper274_U0_fifo_cin_in_V_V_read)
);

(* keep_hierarchy = "yes" *)
fifo_almost_full
#(
  .DATA_WIDTH(32),
  .DEPTH(15),
  .ADDR_WIDTH(6),
  .GRACE_PERIOD(5)
)
fifo_cout_drain_PE_12_2_V_U
(
  .clk(ap_clk),
  .reset(ap_rst_n_inv),
  .if_read_ce(1'b1),
  .if_write_ce(1'b1),
  .if_din(PE_wrapper296_U0_fifo_cout_drain_out_V_din),
  .if_full_n(fifo_cout_drain_PE_12_2_V_full_n),
  .if_write(PE_wrapper296_U0_fifo_cout_drain_out_V_write),
  .if_dout(fifo_cout_drain_PE_12_2_V_dout),
  .if_empty_n(fifo_cout_drain_PE_12_2_V_empty_n),
  .if_read(cout_drain_IO_L1_out_wrapper402_U0_fifo_cout_drain_local_in_V_read)
);

(* keep_hierarchy = "yes" *)
fifo_almost_full
#(
  .DATA_WIDTH(32),
  .DEPTH(6),
  .ADDR_WIDTH(6),
  .GRACE_PERIOD(3)
)
fifo_cout_drain_PE_14_4_V_U
(
  .clk(ap_clk),
  .reset(ap_rst_n_inv),
  .if_read_ce(1'b1),
  .if_write_ce(1'b1),
  .if_din(PE_wrapper322_U0_fifo_cout_drain_out_V_din),
  .if_full_n(fifo_cout_drain_PE_14_4_V_full_n),
  .if_write(PE_wrapper322_U0_fifo_cout_drain_out_V_write),
  .if_dout(fifo_cout_drain_PE_14_4_V_dout),
  .if_empty_n(fifo_cout_drain_PE_14_4_V_empty_n),
  .if_read(cout_drain_IO_L1_out_wrapper432_U0_fifo_cout_drain_local_in_V_read)
);

(* keep_hierarchy = "yes" *)
fifo_almost_full
#(
  .DATA_WIDTH(64),
  .DEPTH(4),
  .ADDR_WIDTH(7),
  .GRACE_PERIOD(3)
)
fifo_cout_drain_cout_drain_IO_L1_out_2_13_V_V_U
(
  .clk(ap_clk),
  .reset(ap_rst_n_inv),
  .if_read_ce(1'b1),
  .if_write_ce(1'b1),
  .if_din(cout_drain_IO_L1_out_wrapper401_U0_fifo_cout_drain_out_V_V_din),
  .if_full_n(fifo_cout_drain_cout_drain_IO_L1_out_2_13_V_V_full_n),
  .if_write(cout_drain_IO_L1_out_wrapper401_U0_fifo_cout_drain_out_V_V_write),
  .if_dout(fifo_cout_drain_cout_drain_IO_L1_out_2_13_V_V_dout),
  .if_empty_n(fifo_cout_drain_cout_drain_IO_L1_out_2_13_V_V_empty_n),
  .if_read(cout_drain_IO_L1_out_wrapper402_U0_fifo_cout_drain_in_V_V_read)
);

(* keep_hierarchy = "yes" *)
fifo_almost_full
#(
  .DATA_WIDTH(32),
  .DEPTH(16),
  .ADDR_WIDTH(6),
  .GRACE_PERIOD(3)
)
fifo_cout_drain_PE_12_4_V_U
(
  .clk(ap_clk),
  .reset(ap_rst_n_inv),
  .if_read_ce(1'b1),
  .if_write_ce(1'b1),
  .if_din(PE_wrapper298_U0_fifo_cout_drain_out_V_din),
  .if_full_n(fifo_cout_drain_PE_12_4_V_full_n),
  .if_write(PE_wrapper298_U0_fifo_cout_drain_out_V_write),
  .if_dout(fifo_cout_drain_PE_12_4_V_dout),
  .if_empty_n(fifo_cout_drain_PE_12_4_V_empty_n),
  .if_read(cout_drain_IO_L1_out_wrapper434_U0_fifo_cout_drain_local_in_V_read)
);

// pipeline ap_start
initial begin
  ap_start_p1 = 1'b0;
  ap_start_p2 = 1'b0;
  ap_start_pipe = 1'b0;
end
always @ (posedge ap_clk) begin
  ap_start_p1 <= ap_start;
  ap_start_p2 <= ap_start_p1;
  ap_start_pipe <= ap_start_p2;
end
assign ap_done = 1'b1;
assign ap_ready = ap_done;
assign ap_idle = ap_done;
// pipeline ap_start
initial begin
  ap_rst_p1 = 1'b0;
  ap_rst_p2 = 1'b0;
  ap_rst_pipe = 1'b0;
  ap_rst_n_p1 = 1'b0;
  ap_rst_n_p2 = 1'b0;
  ap_rst_n_pipe = 1'b0;
end
always @ (posedge ap_clk) begin
  ap_rst_p1 <= ~ap_rst_n;
  ap_rst_p2 <= ap_rst_p1;
  ap_rst_pipe <= ap_rst_p2;
  ap_rst_n_p1 <= ap_rst_n;
  ap_rst_n_p2 <= ap_rst_n_p1;
  ap_rst_n_pipe <= ap_rst_n_p2;
end
endmodule

// first-word fall-through (FWFT) FIFO
// if its capacity > THRESHOLD bits, it uses block RAM, otherwise it will uses
// shift register LUT
module fifo_almost_full #(
  parameter DATA_WIDTH = 32,
  parameter ADDR_WIDTH = 5,
  parameter DEPTH      = 32,
  parameter THRESHOLD  = 18432,
  parameter GRACE_PERIOD = 2
) (
  input wire clk,
  input wire reset,
  // write
  output wire                  if_full_n,
  input  wire                  if_write_ce,
  input  wire                  if_write,
  input  wire [DATA_WIDTH-1:0] if_din,
  // read
  output wire                  if_empty_n,
  input  wire                  if_read_ce,
  input  wire                  if_read,
  output wire [DATA_WIDTH-1:0] if_dout
);
  parameter REAL_DEPTH = GRACE_PERIOD + DEPTH + 4;
  parameter REAL_ADDR_WIDTH  = $clog2(REAL_DEPTH);
generate
  if (DATA_WIDTH * DEPTH > THRESHOLD) begin : bram
    fifo_bram_almost_full #(
      .DATA_WIDTH(DATA_WIDTH),
      .ADDR_WIDTH(REAL_ADDR_WIDTH),
      .DEPTH     (REAL_DEPTH),
      .GRACE_PERIOD(GRACE_PERIOD) /*********/
    ) unit (
      .clk  (clk),
      .reset(reset),
      .if_full_n  (if_full_n),
      .if_write_ce(if_write_ce),
      .if_write   (if_write),
      .if_din     (if_din),
      .if_empty_n(if_empty_n),
      .if_read_ce(if_read_ce),
      .if_read   (if_read),
      .if_dout   (if_dout)
    );
  end else begin : srl
    fifo_srl_almost_full #(
      .DATA_WIDTH(DATA_WIDTH),
      .ADDR_WIDTH(REAL_ADDR_WIDTH),
      .DEPTH     (REAL_DEPTH),
      .GRACE_PERIOD(GRACE_PERIOD) /*********/
    ) unit (
      .clk  (clk),
      .reset(reset),
      .if_full_n  (if_full_n),
      .if_write_ce(if_write_ce),
      .if_write   (if_write),
      .if_din     (if_din),
      .if_empty_n(if_empty_n),
      .if_read_ce(if_read_ce),
      .if_read   (if_read),
      .if_dout   (if_dout)
    );
  end
endgenerate
endmodule  // fifo
/////////////////////////////////////////////////////////////////
module fifo_srl_almost_full (
    clk,
    reset,
    if_empty_n,
    if_read_ce,
    if_read,
    if_dout,
    if_full_n,
    if_write_ce,
    if_write,
    if_din);
parameter MEM_STYLE   = "shiftreg";
parameter DATA_WIDTH  = 32'd32;
parameter ADDR_WIDTH  = 32'd4;
parameter DEPTH       = 5'd16;
/*******************************************/
parameter GRACE_PERIOD = 2;
/*******************************************/
input clk;
input reset;
output if_empty_n;
input if_read_ce;
input if_read;
output[DATA_WIDTH - 1:0] if_dout;
output if_full_n;
input if_write_ce;
input if_write;
input[DATA_WIDTH - 1:0] if_din;
wire[ADDR_WIDTH - 1:0] shiftReg_addr ;
wire[DATA_WIDTH - 1:0] shiftReg_data, shiftReg_q;
wire                     shiftReg_ce;
reg[ADDR_WIDTH:0] mOutPtr = ~{(ADDR_WIDTH+1){1'b0}};
reg internal_empty_n = 0, internal_full_n = 1;
assign if_empty_n = internal_empty_n;
/*******************************************/
// assign if_full_n = internal_full_n;
wire almost_full = mOutPtr >= DEPTH - 1 - GRACE_PERIOD && mOutPtr != ~{ADDR_WIDTH+1{1'b0}};
assign if_full_n = ~almost_full;
/*******************************************/
assign shiftReg_data = if_din;
assign if_dout = shiftReg_q;
always @ (posedge clk) begin
    if (reset == 1'b1)
    begin
        mOutPtr <= ~{ADDR_WIDTH+1{1'b0}};
        internal_empty_n <= 1'b0;
        internal_full_n <= 1'b1;
    end
    else begin
        if (((if_read & if_read_ce) == 1 & internal_empty_n == 1) && 
            ((if_write & if_write_ce) == 0 | internal_full_n == 0))
        begin
            mOutPtr <= mOutPtr - 5'd1;
            if (mOutPtr == 0)
                internal_empty_n <= 1'b0;
            internal_full_n <= 1'b1;
        end 
        else if (((if_read & if_read_ce) == 0 | internal_empty_n == 0) && 
            ((if_write & if_write_ce) == 1 & internal_full_n == 1))
        begin
            mOutPtr <= mOutPtr + 5'd1;
            internal_empty_n <= 1'b1;
            if (mOutPtr == DEPTH - 5'd2)
                internal_full_n <= 1'b0;
        end 
    end
end
assign shiftReg_addr = mOutPtr[ADDR_WIDTH] == 1'b0 ? mOutPtr[ADDR_WIDTH-1:0]:{ADDR_WIDTH{1'b0}};
assign shiftReg_ce = (if_write & if_write_ce) & internal_full_n;
fifo_srl_almost_full_internal 
#(
    .DATA_WIDTH(DATA_WIDTH),
    .ADDR_WIDTH(ADDR_WIDTH),
    .DEPTH(DEPTH))
U_fifo_w32_d16_A_ram (
    .clk(clk),
    .data(shiftReg_data),
    .ce(shiftReg_ce),
    .a(shiftReg_addr),
    .q(shiftReg_q));
endmodule  
module fifo_srl_almost_full_internal (
    clk,
    data,
    ce,
    a,
    q);
parameter DATA_WIDTH = 32'd32;
parameter ADDR_WIDTH = 32'd4;
parameter DEPTH = 5'd16;
input clk;
input [DATA_WIDTH-1:0] data;
input ce;
input [ADDR_WIDTH-1:0] a;
output [DATA_WIDTH-1:0] q;
reg[DATA_WIDTH-1:0] SRL_SIG [0:DEPTH-1];
integer i;
always @ (posedge clk)
    begin
        if (ce)
        begin
            for (i=0;i<DEPTH-1;i=i+1)
                SRL_SIG[i+1] <= SRL_SIG[i];
            SRL_SIG[0] <= data;
        end
    end
assign q = SRL_SIG[a];
endmodule
///////////////////////////////////////////////////////////
// first-word fall-through (FWFT) FIFO using block RAM or URAM (let Vivado choose)
// based on HLS generated code
module fifo_bram_almost_full #(
  parameter MEM_STYLE  = "auto",
  parameter DATA_WIDTH = 32,
  parameter ADDR_WIDTH = 5,
  parameter DEPTH      = 32,
  parameter GRACE_PERIOD = 2
) (
  input wire clk,
  input wire reset,
  // write
  output wire                  if_full_n,
  input  wire                  if_write_ce,
  input  wire                  if_write,
  input  wire [DATA_WIDTH-1:0] if_din,
  // read
  output wire                  if_empty_n,
  input  wire                  if_read_ce,
  input  wire                  if_read,
  output wire [DATA_WIDTH-1:0] if_dout
);
(* ram_style = MEM_STYLE *)
reg  [DATA_WIDTH-1:0] mem[0:DEPTH-1];
reg  [DATA_WIDTH-1:0] q_buf;
reg  [ADDR_WIDTH-1:0] waddr;
reg  [ADDR_WIDTH-1:0] raddr;
wire [ADDR_WIDTH-1:0] wnext;
wire [ADDR_WIDTH-1:0] rnext;
wire                  push;
wire                  pop;
reg  [ADDR_WIDTH-1:0] used;
reg                   full_n;
reg                   empty_n;
reg  [DATA_WIDTH-1:0] q_tmp;
reg                   show_ahead;
reg  [DATA_WIDTH-1:0] dout_buf;
reg                   dout_valid;
localparam DepthM1 = DEPTH[ADDR_WIDTH-1:0] - 1'd1;
/**************************************/
wire almost_full = (used >= DEPTH - 1 - GRACE_PERIOD);
//assign if_full_n  = full_n;
assign if_full_n  = ~almost_full;
/**************************************/
assign if_empty_n = dout_valid;
assign if_dout    = dout_buf;
assign push       = full_n & if_write_ce & if_write;
assign pop        = empty_n & if_read_ce & (~dout_valid | if_read);
assign wnext      = !push              ? waddr              :
                    (waddr == DepthM1) ? {ADDR_WIDTH{1'b0}} : waddr + 1'd1;
assign rnext      = !pop               ? raddr              :
                    (raddr == DepthM1) ? {ADDR_WIDTH{1'b0}} : raddr + 1'd1;
// waddr
always @(posedge clk) begin
  if (reset)
    waddr <= {ADDR_WIDTH{1'b0}};
  else
    waddr <= wnext;
end
// raddr
always @(posedge clk) begin
  if (reset)
    raddr <= {ADDR_WIDTH{1'b0}};
  else
    raddr <= rnext;
end
// used
always @(posedge clk) begin
  if (reset)
    used <= {ADDR_WIDTH{1'b0}};
  else if (push && !pop)
    used <= used + 1'b1;
  else if (!push && pop)
    used <= used - 1'b1;
end
// full_n
always @(posedge clk) begin
  if (reset)
    full_n <= 1'b1;
  else if (push && !pop)
    full_n <= (used != DepthM1);
  else if (!push && pop)
    full_n <= 1'b1;
end
// empty_n
always @(posedge clk) begin
  if (reset)
    empty_n <= 1'b0;
  else if (push && !pop)
    empty_n <= 1'b1;
  else if (!push && pop)
    empty_n <= (used != {{(ADDR_WIDTH-1){1'b0}},1'b1});
end
// mem
always @(posedge clk) begin
  if (push)
    mem[waddr] <= if_din;
end
// q_buf
always @(posedge clk) begin
  q_buf <= mem[rnext];
end
// q_tmp
always @(posedge clk) begin
  if (reset)
    q_tmp <= {DATA_WIDTH{1'b0}};
  else if (push)
    q_tmp <= if_din;
end
// show_ahead
always @(posedge clk) begin
  if (reset)
    show_ahead <= 1'b0;
  else if (push && used == {{(ADDR_WIDTH-1){1'b0}},pop})
    show_ahead <= 1'b1;
  else
    show_ahead <= 1'b0;
end
// dout_buf
always @(posedge clk) begin
  if (reset)
    dout_buf <= {DATA_WIDTH{1'b0}};
  else if (pop)
    dout_buf <= show_ahead? q_tmp : q_buf;
end
// dout_valid
always @(posedge clk) begin
  if (reset)
    dout_valid <= 1'b0;
  else if (pop)
    dout_valid <= 1'b1;
  else if (if_read_ce & if_read)
    dout_valid <= 1'b0;
end
endmodule  // fifo_bram

